// Copyright (C) 2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std
// ALTERA_TIMESTAMP:Thu Sep 13 06:32:39 PDT 2018
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
iNpb08z89KrKBdR1cAeEBR2lBFqkgkhYP8wPfMabYFfzOigkXG0OAqK0lgiJTlDg
zl9ksH9Ndsb4QU3/KU3PuubMWQNWUmytYPX5aBP5YNuLBi8xmPEceFn926seakOx
Y0/5FMzBYJnv0OI1Fer5ZWw8txK5j5YtvfwZeBWOSyM=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 28208)
X0Zm/a7C0Fyhd4PJHUAIR58xAel4V2+LttDtrkTvRC2Ymvvh/sGeHFGKU6Fjo0c/
iSsSyZO/7qMecZTpFiXkYBvLpMIFnpYPxxInCRApePPDq9Auu/UkQ43/w98EYGpr
KNGFabExbvLrMSbYJ7VR5/LF4ntuU9GaiwIDLVymSGxjM/ebZWdHg63jfU/WEb/F
JYJ9ZFN5EpIYAQ6wkPiSA10Kea50UeiYKhgcYfE6HgdLldJd94WWSBmrYOzk1bPA
1UF84N6gygY6xHftvkM14WvwJ1vY/RzbJrXJFIlObtTfqMVm3FD5oZxisDUOf0uk
rXzXNAF5LmJwOE+MmyW3DTKG/saQ7nzv2o9qRryTq1lDsSEXJUwMUuLazC4/xBnI
Pi9r0uFZgbaGOfI1/uvyRjFfKzLkWYO/QNVOj6L62aEz0MAzIqqtfAVhx+CtsgpC
RMRISS//rLBxhig2zgKqZGHUzVwrPCdpbrwC3536hE/jZq+QrFuyY4g7Y9/EvNZ7
rmyH5e55hvtgSX2DvxxHdZDrP+MWjIwh43mhrsqRWt0gcsRAIZPNaXAYwduho2AE
IjVSFhzWMDptIEmeZyOGGtS9Z9RBCAkJ8atIoybwcueCmVnDF9VjcGM3WFgm7eNq
FMCcc3zgbs29G0n3iJLBkUMCdmJn5zZgTuN0r4gQxHzE2+Aq1U41SGXrEOOAoVeE
ATVjHpK73B9enQ7RDGLcOdZ35MEZCPmLFoWu4x31v1wdkmX4tOfccwJkajgTA7rC
PnCHkdTZVap1rSYpsct9q2XTLvbbdWcr5BygHramd1/V5LdHOPmE8Jpz+SoKNI9a
gXcdbjUzqEZkrhBket8BruVUYyr1zUp4vgmFz+fK5pN0xTg7m70cyx54R6UwEihE
GgsOdIiU22RNa9xC8ozSozoIGIDbaE4n0dykW83b2Hk1tdB7cq/U//zsdmKgF93c
QkJA/vef6gU200XqqNeRX6gqWiwZxFyjKL47yBhHA7CerbTQBwHK4CfaO/9Lp2gZ
nIgPH/kkTHXVYjd/KRosgdep5RajOE1tIYu5BsxUXuThL0jAkIM8DbwouUkCr7Gj
EaYHZ3v+f8fygLtJgr/Ziwowu3yfk2tCk8P6auirVJnlzPb5WrbpagKrAl/P4HMx
IbULFL2Hp4vrsGroxl29aoouzz7Hdu+yQfNdREIIGd5Niux6uML3pnXOx/8NRanx
/7D+sk0xcO6RGv25e44Xq10ps4l9QL9EBO/YNJ3mvvz2wqZNfSfA6xmyoxMhuAgb
1gVLDv3gBzEPxWzNMJnyUk6dUwZwvlWUOfoDah/5er6QAfUcQ7X0opwst+nUaLbn
YkzokrTh6+H2PJSnB/Bu1wpCbs4Q6CdRBzmXDYm/VDa8hihFgZr5FUHn+GGVe39p
PVIRdQF/AT8fkL+q7vd9+teAUXK7UvO3oJcOgmcLS2Z1lB8Dcqn4fQEdp4xBkuMF
dSYcFmKRyYZf2JSe6Sz0qqJUdliVq1RzMLssEKFYsvpSlpaPavUhY1K8guMCkUm/
HW3acLRmY3/IuHUwjPAZxgaMrp4vu6SsCYSyadDuBjTQjteBD1665fXCjPq6wW4b
tEIAbj3g3rPbY97xFJsOVsbGEPKAdVQlfZb1+/Acx5YmwWIXGJ8w1tZC/R9L/NLq
6Le1AjUJAc/17ZtxF4DN6UsGqulxcGMh2QG3HVdwMXcaM4cRtvxOSX2JB+bLA7oZ
Rjg2AMIfBNI2qOAL/qh2NssrdWvkgTHbWGwgNUazAwmvS7itWsvzVz0l/dmHiwoa
UhQoMdBhuaoA0gKAubqlI8JstuA0hC3mnYHOz8m/soLfSi5AIEDUc3DXXmo225ec
2tTmMMPK02dlWcOwbp5tgPytSBBUequA5p3IC1P24bffc8hwMFNPPomVf5BvvmwH
FhZPc4dtNF7C8OO7PA0q+OCHHqhmL85ZsILM8lpTC1BoW7en1eCBqMLUauoERHpY
XERDP1Oi38ou+LJaBXXbj2a5IKYvbsddQSJywkBXiH8Vsc5lvDvK5FYHxDcwhCva
tjx8kHI2TysYLIvDnaPJ7SPSwmj5/EFGD38qmO/nP7Lw0YHbiDczG0soCAxjTXQ8
zTTCwZqMM12tHw6lBrtgsZ60ukGXfpd9Nwqf65ZfV6EECIJS+b3w4hT4M8Iw2k2I
0DL8gq7O78kvRp1qllX+tmUGyDZ4AlG5K13aXRNhQlfMx4QjckPkh9HEM46tl15+
d17n4x/HXucIpVtyz43AVqcMA8hmsTF1VZj8EgMVz3eg1M/mM7M4YcQOG6swki1i
hdUVkZPj+VSN1JMZ427KSdLP6D5J2XWL3r7NvsHKrLNoxIgtj4u2U2zBrNuWaoRU
c3SAjzy+if2mc8drSLMC75nKq7dTiNnE4UxksTW6Rg1KoAsRdj3lluTEz3xaLEDK
XwqtDFhYUgWl0Hqj2xe2NbIP2ipd/T68tSj45EfxcvQ4qDiicpqlfC0/6UqPFdPg
ukowbHZl5NdMi4myKnN4Gs5bMWfrdQji/1Y0ebBlhpkck3xMX/E/jddx6VvDhUt0
ArB5Zc+AE9jJVkQv6Vlg5G3Kvf8Zy+9ZezXQhDBQaBc8JJa/K1RwLL68RhLb0it0
Ob1e8aDkDXVRPd9C/RfUIv1XTlSJqYH1JSAUGfZ6nv5KiVWUYzjerkrFVPKqhBXy
bbO42udF+kPTTMHnHSN/QyJlea8SaroMhp1P05FN36H05RqApNYKwLyjGsCR9vO/
0UhnJEwL5OJy5yVs0n8YlGR+JXvPiDWDp0fyZMc/EmNPYY/VBKLXFs2KLTKCzN8M
8BLLevMIW4QAka14uwHF3l6ejcTKkc7uvQDbnIXdf8tTHJYfTQbrvAbW3hHVUh/R
TGQ5Jl0wph217ndSAkr7Ob+LSvoyehbrjoTlVAsEd++Pbw9+4922rATASsg9e0nL
sxTvoWuEhtGNdpvqTv3a1YaJlzOTeJq8HPCjl3lFtzF664UcDT/NoC+7JYDPkTJP
BFtYuWLSQ9Zt04dVXSsUCNKuSrXxCz2zXm1nUWuSLP4c+aSgWh2Go3sxm2VHDHd5
pj5I6yHzC0AdiUSuBEf4K771Vu6jr04Blue7Sa+Ga4eMRowK6R5JN3144G45dWG0
Gmmq+5N/TQ9FihVjy+k21YbFb97OpD6OvzEb8KWbOcQwJ8KTFrB+V/9mPipF7eoj
JwYXlqWbgmePvYb6RiLihAQUrV9FDx/3SJxvXqK3n13VtbfnchcYGGXj+YzQmAoO
oWB5m25mYNdGN6G8mr8fblNr7MX83zhIHsuN7nikyfdW9TDEJC1hk4DMe5iUeoX9
Pj7wLfcl7bGNmum1w5FWRoUHHGAs8+3BFo6HAAU/4ANo3OTPsNMGy1NcfJTHgTXP
Ny8P9oHHNx9t8jvRoMUJr8uDmCzinl4r/zMN0aKBCA3avmeUN1Lb2xV2Yi7N2GfH
j4mrSt15psCGVO1on0+zTg2QvuvjKbXmG2taC0ONvXqoW2hWdZu+nJslRScnizSa
ogSIWAQEKl9XkSo8YbM9mYQtehJqObxLA1d23atG79Wu1l5pJU50kc+gUI4G7UTU
KArjk/vtA+fKYyEf8LvailqBxAAkqIYVGJ7b53PA7WKa/0youues44Zn2Juu6AUN
ZRH+CRjOEb6vyLksMV2BxftXt8yNaueUUX64hrXsMbDd3XPYA4+2o/3tjlOMqzeM
JecrrS7dlpBw+40WCOb+y3pgNbTKr3ISj7bpUSn+vikBJGxpa++uCMf1bKmw5GZz
P9IUy5xK+qpUxWOekUxdP8HfEBvfKV2dbsRa8/vwqiCC/hjaD9FsGq2fapD/29vI
RCzhdPIeRX8pwYHRVBWu+mroySxA7uaAb9XvOAwxUztufeIoZPBwA9AlKyBuFSw7
t3Olt/r6pA0+8j2ZkkVNxI2gyGYiDaspr8wmKlU7RDxNP4QBHmZQPfiWBVdXkwmg
iCjI0+IrGlYCS5sa9B2vJQUxPciMsn4gcqSkZnfrp2Lpps+zKT4/9szVra/Uyhcd
a4FnPREFp4MRls/KWrp0WHUpGCB/xtfTqK8s7fgBpR+1mS/+jS22OoGS3z+0rE2K
mtiJx7qzRORHH/+FVxDkmaX1xzE1m27CN8jOgyahYMQ1jxwgH4o+SHQIfeycG7fw
CEkKfkoPmXDpm9XNTqxS/Yxl0R3MnM1M+uAmiz+b5Ob4k4vbY3mRt+blM9QlvYuz
Xgy6ZmKnV4jhlITAcVMbu/L96j8Tf3ADDSgSmSepQgeNz4dNdaSLr+c090lA/F2S
LH/QTaU+XSoyfD+x6Tr/0ZqQI5jEl+QUzxx354d3QK6E+U4qXjuL9aTDNKaIAIYF
WYRigdUnoywrQUdOANLembHy4qvLrlqV0HPBRbacvGPLL1PpvtxJPMjsb/z+4ErG
huhrWUsbob2eZ1SVYmPLNqdV1i1KSXiT+/JsOv0t6Q3/11+PyuIiXEThIc0+HURa
Dd7rAw4RYru1YegF3crKrY1ePFU5Bb14CbHgcF7wzJi/0/wqHDL3mQUQHibyYK0W
3OvEZBjTeq1tdzlohfwuqABrIkGwHDfMi3UkrmH7cvpmN6dHdeL5JcCDieBTpWA5
Gf7qSyT/VFWaKYiGv59eCucDfJeuJfKbTY/2x1MKcvu7jqHP2Yn+wmyYNOxXvz/z
sAkEDRs2GhjPL4wWWRlXh7c7wytbOIhpMzSufR1sBqKBZFAyagP2Sy3yDKbc+xKZ
qV6yj/vbgFAuQxnMRVbTza0mC9QFW6dmsojHc6LI6S2f9bcTcjMJDN2nw5RCwWNJ
WfZ91259XV91I+F+fdvBV47BnFARhTXibbfQIvwD5i7JbrZFFBHQfcP87Rdhx0w2
V73eBE5DPEQyPnjWfhSpTPsyxQDwYM78pViMg1caNxO9MeEroWp/YJ5+V3XM90AZ
zT/R4nzgg+kPQpDJxiJs+eiCGHLaVYfCaTjuKoov5n4J+/Np+fFgpfzBnRrNurjh
87kZMnF5M4zlPCOFIGzq5z2w6eDVJfpvEk2l33IFA+wMIKVRkMHaoXANBYdofrWn
S6fajVzO1e46g9SKbQPvBst1hrDZg/kNgmg9YeY+y2aPHuOx/EHWwHBJfM7PUwoH
/9i110KrR9NSr3zNXrE3lHrv3DRg3s0scnw7lr76pI4AmSNGpWaWncV4tOwWGFMV
CuO580IHvj5+qxezCurTRMWjcoW3hUFceFNNq352q9R4OIJT29mEz+ff1IfHCYuk
7c2yIllTOmeLvD+fRSj9R1fF5Nfj8ktrzxWjisk0OFAVFuFyfbECEZl6FrUikh1Y
KWyQbuVKVwP/cCzMpdU/pyVzM/por5Xjgl5lk0VIlFEP99pmGCAJXMtJPQSkGkIy
KPJehzD2q6EDl+tTXHtUhBahJyeJMkuorToTPtdXEcT7Rm3R+okIbdU/a4niKqk+
Gjvikg2AjhZNJSympxz3X/QP9lKzx9Sou7/CLlAP171mA2WHrZoMeziPZVjY46gE
Gs/KwkYc+85cKzPjKbZXaz7Q3E7Wq6MB0qvC0E0iidxGUNjCTNJrkEisQ03H9PGK
ZJnq20eoI1VrNMzJfwGLRPyJqnumbeHO9ZVLR41hfxRvh3q+Xc9L1gDxEPoblXf1
r+OXdR1sOW3oUL3y996BSRwhiWTq5hv9taTVC3cRc7J6vXTw9OFD89nrA/rKKfK/
rf99A/1Tl8ARrdhybL2x7K96YpEz0035jGnuZGASYFXLCTcZPK6RGsiIh40EnE0L
urL9CN97dqBrEcbpKlTAc4QDKsArSiR8LszGBYAwiP8858xJSuyMrdqeZuIEM7vW
Z5kzIekh5OUzvqEBOi5UzVRCzgsRYG+HG+jYWbOLcOzrnO5K2R3Ax8zJNwlIoOBk
fL76OPkzO5dO08bOwd3ZYqZwzNlmXhNZQPgF+os2bjoZ3iykjfJaXBqHJ9NsaF5Y
34JqzHdAnekSxvGQiU+Bme7ZpAQ+yRMiq9ys6FB9dBxC67lVgOXrHEx9xna/W+Cv
ayQHDnq++h77y88Iee2BCeH9dbOoK/TyMQOFDiriQFCwFiRVkqlMwUwSNLX5mNQU
ug0PjR34J3WeOAJKUzLyCqxv/Sha9xVVIZ5kWzU1M1Vp7De8gZPsTuMAss1Jo0Dp
yzpYXDhogXK9uL/lPxjupwkshsp6ufHduyH5iieu/Pn2g9sFunHKnfDF0lDIh+U9
MWiAl37SvewN6y48xGTY4mJvFNmFALVOEuyktQkab3xicCzyHVpPgK+ilLimzhtI
dSqqhD9zdSPxhH0mEFbgoKL1+FCO5rZglt7QypImpKSWTg/DRIMvqJECCvqHmgDD
R/syjnZ2A69bHy9uHIGJrMPPbBFkkJWF0licko7jj4Wurs2IhVQEBNLLv7nvY3yO
oU0y0WZxe3LAfVweKPrnsDjYjtMhcct6s8McNy74fx/BRBVEtjutUalVOsU+CA3s
HpGJKGEdF6CC4xFLhlDIesMXg96MYjG/CWDTxXhQpNJKFs9XVEdHdY2e6D027mYU
jXjxhCsXIGvzGmF/p0TC736Tmc9T+d5ErWNlQobaFw2oubgVBVXRW+CgrBxJIp3t
jBdSAFK+sPP1+9jM6n/FY/oTMj6xFd3YuLbZCYYkPoTNzKcrb+qgHyXDzO+8xYlu
s0Zvf5Xl9Bfy1l6WWhuhOzulXy+FwcgRHA9xiZEqnJxh8XCOxmeEhTFi38C6ZUj2
hzqqWNd+xE3oVWeRQ+/uHIgQS2yGma9Rsd0qCD9XHZ3C8R2p2vVd1b4Uir7LcsMr
deztlmsFAQ0ka71l2DZEK53RZJkR7CYhxMI48fkx39I4nUIWte8dTO2N+OkppfIF
5du8SL5ifk9bdY1dgyZYRyl5Ya9p4Fb0ZrKcttI7W/o1WXFrMNTZHBf8vyE4d9BE
Zlae+W1n9LkYXLzScNBvqJUPvFdVmBVcPIwxAlBjdI9NukKEnP0P2T8MicwiwD7+
drRClp3U/IFSZ1tc7o02zflGP7ZWJnQoKHkyedeqQdJkHwUWAXqGhCaENKQVlATh
W7/K/ChAhTEBV39ADEFfW5YWB3npCM5/xaWLwJR2C5F8BNxUzM2wT1VWuTo3CuZt
AofMl20IGkPdM+PWcaQOXYPdzgYYilv5B7DA/bU7TzFjL2G7O6x3Kt1QNjq+HblG
lNhptauTjvdmbVVVntuiXXF5ACKz1hqfXVQDMg3hxcwm73AlU9csr0CQkSADHoq8
itoeknMCxH6gtib6GiVj4nxW4IeQ2hAmom3MLVh+70DICSH8zE0Q3WPxdzZs4vOP
7Em3ihNcqo3T11HlLXV6mbutvyQJ485Z6DHsq6B1ydBAHQE+DjPqPghwU/VBjYwX
w8RwspB0ES3I74HJXe7Eaqf5DqzcY6L6HNj4sfTyWayNo7c1oQDMwjFhLdD6BoCy
o09fMfRla5ZnhmqCKv6mJt5oS6LaG3HXpRkcW+S5rV0MT7YCKINuilnQ8fdxKr4U
6uuHesKv3ubRW/FcdgCUmu2RvVsFIAwT1NtWgGqFuyuqvHsfk/JtEVf3NRbm/rj/
vO46EAUMGpl84BpcrVLli8BrUw2gBWTasuOHlpepDK2e50q6QTq8jkjnshjn7hIX
vUJTvSTmawrbwSgvRoMM9CsZGonx9Q4y0Zac+2X7w3WFXKgzUzwLRNZ58gvNrIYP
8SlVwqsw9ScBWH9xGCZS+S2DCAdagOD8GvXrgKa8N1/m7sDnkghFXJHoeBqT80wd
TPf1uZBEarXbA8yoOYib74IxmJEtB0q/xUU47J48rAFT6RVEqkgcpI3ejUSfPYXj
cdEr9tSNvYPEv4d9C7TkXLKpT3jNGX3UOuQnPqXvzGg/rv2ysdDwO7ErK/OL5xET
62Nje9KD2b9YjGid5wKrGDnVI6yYwdABS6SmLMeYKbjk+DJSTkJUuMDNNbCoX+Oc
JRYtNhBPErkX7SjAeo8J1j6+qxclFY+g98V+JmAlc3pf3LzSlEH+UakbMSMyF8jL
6o5i8MgLTYGtlMh1J7U+L/v+t7E+e7fULK41IfTtueWJzFtBO0MKJ6XFpz8xpMFt
WC4rRzzOXwWJ/ecKSXfO0wzZvm38XLDoDS6eRc9ISRGpBTuYPYKovjtjhB/o4Qji
KIhLZcWt/3m6qvGjKzdSFH02xqimNxYkvBNDVOgJIuNxVBneDGgR3Irdcxf88GPv
b230pkortjqhqI9frbCO2XHGmskZn2cJsP+1L4urULRAIf5LlKlt/2qtse6hoIYy
RKbzpnrRfd4HCxY9ojrGADe7kTpWi3SWoqpa7KBoBY5Bgzb+UtMMmKwx+oA98vy3
RuoM4YwppJBgfxcwf5l2qKb4LKYkI8bAErDbbfO1+Jy0hn69m3nYB19rYhu2F7x4
XTD8dvEdiA/HX2bfjfwfjjf08ARMQemUNZJtjj4DJxF9ezD0nF4kt3U4vqRpMIwV
kVhdTUwHK6sXEZR3xNpzVMK0Bg61Rw1G/x8gd/xZDAmQzyImS2R2xotlMBoI9+aS
7v7XiLTnq3mck4cvVS6Wvt/EVvLXGMpPJTjKuSDKcyo36em82JxUESLi99Fy7j1X
xmP01hdr1yNe3M9UenVfM5aOfC5qpZttXIsUsVsu56qks8BiC5V145HPDRCbFva+
omTn42LOt4QiVjZIwJ9wFzftoLaA64zXw4oVYkKiYowpPlfccQSKpFP06/m0j1ec
Lzp8U2Tmu9v+i345ofy2rkWawpo6sPLcxeCFdVPNa8lJSUVlfdG8pD7KQfZ9drcF
Y7NFVlrwaigXZYx4BMt1gJ3tyCppVjXup/KAIuw3lV/V37iLoUG1oBGFQlwjJIWC
Wq8y9QtChC5vbpPrU+O6BQVzpsAz5VYZ5HBmWo4InmdmyI6Kv+Sa0znR9pMduXwX
g2CFk1YtxUJSptNAJ1SfCzjdQ8y+bpmq9dmXIL88ceY7vJCMOziXdjrQK2RdJASp
S/I6foQf4vMQSdCUMWuWtg0afKqusq3St0EXjE2WjkJvr9vC1lXhcidKkbta28ws
zg8AzZZeQaboCFwwDjT31i4DQiI7V21SZt/8JtH40Rl2CslHf9cMsVedLtmQ+mfB
EumiB2YC1V6Fs9Lk3HPFb3BQFJ1t6nshMZN18wygz+j9QX0qVeonvxNg+dUx52A0
5QZS+sJzxMy4o1F+BQj4avjMWFzyhluhWTOGUgnBG8kj2SKQYuKoLkds2kGDRjTC
suXsnLSEQQh4Cb+dzFin+3f3BD9/4A5a85H+FpW0ZhiNGE1jkDAgCOl8i4TpsZvQ
0L+4UTKlMzWTLXK2nl5hT8OEKZDRT5SdIaeAWZq4/aBlTmHt/F+6j2kqoaw8pTS5
cvbLJjRfMiraJN6OJF/8NUNYIVMY9osqrIipn+3CUV6QdGNWBApdtHDqc1NmAGqH
R+ZOvriEAEvdRJ0EjXKgq3EKvk+5Tz1QxmiyfukPWHwUHsv6VE7pkWEjhtWJLnlJ
6eIkjSTdA2vnOaUjpFR0+muKRC4e9kM2szwiviR6W6+0/m0UJDN78bP1Kno6IyOA
MhSUJHva9KW805UZAhnCwcsLxopBQJt44C0wmvk1UuzrSF2up5Bfe40YpbWEueru
m12HCbdEfNXspBiMRHFBDt2agF3bk8W3e/fjdESVwIUtX4qyraL/5z/SnrmTQJmr
WbWR6UTZGPO7J7RBH5AyfWIBRFnHR5LQjsSPk1oqaqmDLBMpgb1LZgOAWPC5tI27
KPEBmF5KhlXUIw+5HHDcPLpklfVGtHUdLqq7g0BWZtpXdQ27MfeC9J3apzSMSs4j
0x9mj17u13dt3nmJ/CirhZuqcrA8vunbTiM2ZHNI2/6i+kNFnIjPw1Iokck5Lb1v
h2LgkaIk1KRdbTtxshSyuOK18FGtlBxEhbcorbbpeXCghxkoseVhLQlXvr5AVOPt
Q1PyLIDo+/uL0CBiAoRoZYytl7mNmD3M/0Osqx5vLUBM6uXdJ411xv9f3HpLYb+V
WnCMNSUq5HTafOUJF8rxK65ETZ4/9xMloGIWoqpxZ5xaJVe9l1cPQ/TCzU0FQIWk
JwSHZRGM+ES8iLg2rS0oZXNnFu6Go+VlnhGGQP2ww4kNAbgISMzDvRoCfiGzScir
1cAM2PgfF5HMqqJofMIurSWZ3Noah/efHaoRtWgeIdA3tiOvGbrOr7md4O+1fQ/C
7L2qtwgVXfFYaQo/uI4vrTPRNggwYtX/G63NU+8x3VVHa3bhK4WDTC/gV7/wp9qy
Gkbp+halQ9Uwg9GaqUettp7rb5md/AcuhQlX7z2BNIiiBAY/386/Pp5umoh8GJaF
gj9oXyMclGX/pS9+vKkdZm9iBJJzWcSB1f2rfoZoJ5SLScJtcXyuXpCDJjYmcYbK
/CEK5935z1s+7fpLQYAsTXCe9iS7ptC1+eTtetFaS22ULgJ9qFroYQcotSNP1/Pl
w5Eq+Z6Z7MYpN+gCsQFSkNmPtJRQF3jySKV7enVukehpuboEEPyAdcdmlmaTFrlT
EGkYl87zvBx8im+ILwT+Q5KsMp5TwiIaBJW7/46CQlOp0ZvJy4EAxp530dIDJdzF
RGun2j+j0B+pn1CTtleutderjGVYNeLhH188FkkK53bgEkBWmCsEiR1IYnz0KYwl
XGqxyksvCnUOu/2KE+RNJqV2gg8mY3UAusmnk6kZ5VMvVSQU2ACLHE5Xk/GZ+8JJ
MToVSUZATeJD4B6B6PMWw+tWX+Ctb97ftlnaJ2Pv50ZYpXwzZp8so2LOonuCKD8+
AF7XRN5dXHkf3r74ciuAlwIfWb5l7M9/6VBBFTqV2rRwgRHzvA7U5+lRcOxcdOux
32pql5/ZbE9qeYRk9ChrrO/9ob2mXs8tlhaAq5ZJYVFE3D6OpSaukNDZtoRtq7dT
w3oq5dAEtKcYR/Kzw2YIZmPyB292C3X+KYkL6Q6UdJ6SzN/QMeHDE+mBBdDW8dqf
5OHJQK+0LaTZRE1ynuH+q3F4jYkCvvhZlSofIg96PRaJrVVcr9nsrHRxjVv8WtV5
JT8ihKV84lH7yP/095l/WrRtaxmCLMHnF/+4EY0DHcMaSJZl1AY1l+FnZuGoRv4q
imcudr8Hcz4VJcjEmgx4Nrn6Ae/6bMB9L+3nygnJ9DOu8aT+8DbsX/pJSz1qcTv9
+hCr9PUW4kcY2qUxNs2v66Rhtei4r9zViJste4KnvNWvqEpaURq+VquES6OzSSWu
DaPPbynyA8D82wE5+rU/bc61YRZYHWoFq2WoD8BQmyPCKnJNopRDqxpcg6JzZUc3
1y040aK1Yf51HRGG8GQxAKl2WjY3Pohzkl5RKbHNzjpjO4ORyU7aYtU9RZjv5CuH
bRaWYSm6UDsrAzsxTs6UIdLPePSY9HRwHKfV74mI+B5RXXdiensjRwr6ZWgY9Xkt
amuSjJNqGclLiQPnK/H1QF4Fngs8eH8xliGlRFH5wcs7bR5sBdEbmloWXnQ0qsZU
avw12GBfnO0qjFZzFd7cwC22kJ2/aS1NiQBL81xVOVf8r7q8Nzo/fBS3PWdFor3Y
QuyTRxoGzV2Dq1PLj0T+sy+CINErX6r7HkO/UcUIU+50/mEY/8SVU5O3dCtGCGFE
lp4shOHMsRUsiwvNPfdY56k7vfUrJjj2B5XFw+y/Pa5p7sm9rOJ5Vdl/CT3rQgMT
Bp9G+CBrWPcY/BeqdxNdP+L8mbs1G8i19QA0kRrOeVASb/G6CvBsEH4XfIiPEIdc
7iek0inKCLVMuFBw0p9RJq+6bcy0jrVHOJY2DvaOv94dSGuaGKOepHN8/bWun+DV
CjXPn+6ayblA2cvUUlN4d/UnHkA2PAHsLTHqk7bvJcEeBxCDal8OxIITMnfZoEJ1
kbWXBLPrAnzeoskZghT6OQwtVKQxgNuoNcQhxkYfMD3gShMde2C51E8s7lDWuB2j
+bWCcShe6JXtP/kamAiW3AcuYs7Nlo8+3ilL02EAY9TOHHnlLqQbo86z56cgFzes
MqohP8ZFLK4RE1QKaBwIIxY2Z+SWyCMdtu8WueC48eAut04u/tsRyQ3h+6hpsvp5
eiBukO072ZrTpSjdG2l2ehhLD3ECzwp9QxY/aCfIDp7nEZSkR9hQ0jQtm0GXdvqw
gLS7Xd/GskpPhWp29FzaYF5qkqY1m7uXpI+LyyIg2aVIlJ9YoUStcx4RFQ9/dxYU
TInJTBqgCQURaujVi1HkaK/Bvwg4Thn1G9ZBcXNXKSDcObGp8qm545Ivzq3QHua6
GgmDM8YekjCfne0EghpcjyLav13Wd49AslpDhl5DpcPIirGBzMhDi4XXneX5IgKS
jdX9u1mejPDJUOUbBd5nIFH04Ve4sZOuz1NdmifiLJsGARt9FojlbRSZKLeprU3z
J70FhJPRPz7MQOyk4Sk2heoZ6xgEGSiCsqFy4aKGRqgwCHjndTN4u8N0atLR6Ah7
uIffKBUiL1VgKgiqbK8TLpSDvnwRM1L6Ddxjze1Lq/mAdan27ZDDmyr08jkPcV5v
Mj9tTH4xfQ9paEeJG0+wZFzBMkPACnRQ3+D3iV92Zp2FFUzjeaXF+DQbWzSUBaSb
9tKXO/tQROfiS+G3DiwuwaN+55bskVZvOlt46Wc7H+Cv7jRYPtN/VIy7iE38zQsm
3RNe1JSSJDmd8PYMX2GKPCYory8XCFCqfqPwdYiTxGbSZ9LG0KcqnGeAJRfrP6Zs
yMI17Dte3DPCchXSBAaXT4DWrlymYlzYZVaXD+8K50D1foK8xLfl3ycdaZo0RqjF
Rqf2XA9dpRNY/SuCafDnsS215cykyB7ujtlFRTW4DXmhV7nw1u2oUuneB+LEtgWi
6yoIziYCRHz0inzEm1o6m70SpRUvtRKBURM95WaVSAht17zGFbdmUDQmGdRHOAeP
TiFbSPIrd3JquXKLwGPOsfNEgHi6JKFcgHUGX8sV47oXNfLO6ANZ+DbpUgWRtL7R
xfEVYeDy0mK79+hCRUFoIxmasgKCi/ikKzyHcZV6IsKcMTw1s0WjXRmW47Fi96Re
qyLxLzwoE8o6+mIj7liLK0tDRMe0SUyLK7cVFs3chD1g27nRMzFybUDcfiHAa/xj
9XW01+fqOVDQbSBw7Oaf1eP5ibYODx1PlaKbcePg6tSNmOu0GEmMMUhLUXOitxDe
3xD7rBs52dPsR+nDYlIn9MD0OtI6koQ5OQHvU5YhksnYTlpB5lEobHfXvWE/gaJB
ikXuKyg7k2DnnUM3NgEATwj8DNyd+EITGfrGooEnXOs4wuFO1IkwzGI6eKNFiT2m
sVfkXBH+dKq0eQdWKo1MGb8Bc+aeue6fQyVXpm79fouGvnnp9nuVPq/kMaEO+cMN
aMmzgQCuMxJ+gWuDdNy/4RvcBsH/PNEVNnhFEO6IBrezuqQcxSb7sW85OlxHY+hA
nKEROj8YZYlOXOIyHKtnrBuHgalUF/S1nnayJroJwh7Jhvl1utKkEB7KQhdaV2jn
0ips7/si6JkF04Amc2Ct1YeFcikPe2icDNEYzRV6UKXXo5Fk5Te2/7eCcaJJTdFB
XeAQVPK7SqUjdXh89ADQSpxKsucBVdK33YA9CK5zJE2ODZTRzj4p9awfo0gNTSR2
GZ6/hupNNTpGmrjHncOJc/NNuPgHhmJEthZOzqO1Do3V6bORFjoX8rdKPPJ1+E/J
d8yUAt9f7fSZcdQ+V886EF6BYRHfUEI+QIY6Jjte29SKJpzWjr0RptIAk9oBkOTX
giwd+z7mok3WrLFT2lEx3xWvXavpWWBfbita3USuKkumILGW7jwPi65D94sr3XRD
3MJR+KsIlVkmEKet6SjIoAPLK17PZ5iUqgcBMDhOuFjtW4GXtF7HTS9Y/IiJe0Gs
nbfylVhq8fagYAKIrkEOV/TDvGSyccqJJK3SYTiPGWYjYumENVhIJ8m3ECFfF9Kx
OukOHxuVjnz9bxDTciLXZDsHpsecY4uH+fdmyBTSGv+wNpvu/TSLxSm3Z67yugFJ
fOLd9LfoK8Gqj3QJvXuI+49NZf9rUIDYosJ1caF557ffExRdtIvnCsemkl0vqpG+
NXoTpEbcjPGdMGKRpXb1NNdBb8JKj3Sy7wIpAd33IWKY3iIouWgnYUdxaExy7syn
fr6xvHMnZxeO8S/vCuK5JRcgaEdkkfv5VzDhydN0mZbogBC6anzsq5xBai52Jkpx
zd7jV++Mmz3/v7efSR36k6aFCMQt3S6axkr5fbwqZJ6QRvkpu1A2khLHNW2Iav7a
BUh7atfCHIJOGQ6To9u7HaBAVDZnA9Jp60yJwh8Ax32CLO2Ri6plEuwQcIxZQYxw
D2/2X+1KKtxugxpD1o63P6c/lP8O6cuV5FCqvTr7q/r87uTdYsSWtLCdhs5v1P5t
V5yiF2jQxpsIt14Ouebuoi1duoie7qFnCAlgTgfoWSqOXsKGx6ovimy5puuCMMFZ
3AeBRc4noHIhXef9aUhsls9DAAJ8KxghsdvKvzGhHFqWlNKs80xcMdg/r6xXsiw9
57cNRJFTp/33LDKHZd9QiLjKle0Ch1bb/rWLSdC6zKnJSnLrs2KwG9m1dMqIrKJS
IB+rFDMzUTkoqqFkZyV4d0gs54i7HjlLCl/Pl1de/yUnfLUFJBkuQuCZ1UHtOE8O
BKbNLQlDghooj0g3UGJEjuznnrOfTNYXL4YIg82/qkvgPqmaameEvcNnqNrLR691
sngrQhSJiX1BMAhAp2lcEA3pTvMt1qC10dLeyeHDQRhUV3MnvJKblTUD0gsbKUox
50u3jz6l6WTFdhCII38n9CmeDW931NbCTdiDveM3vnOlIfkZle5a/nZ1dmOIo2Cn
tV7afoTBmnmIKAsCOgYbHffcwEYLtppO/jB2AKN+BDCWCvNCeNNeDGlWXIL1BOQ5
BvVjSJ36NGTnCPvkdWAQQ4miI/IzGNIQtGKx1ay1WnCAFbW1bY3TPKe/DAEXbuPm
trWN2Zaz/bbW0cy/pfW121CfwWixpxtft0jiJyhWQw4ETBPrlb1mWTOX1Hl8bIqw
EmzRHpGc2ypM61OZ2H4J5UmNihBdcIQPY+LHZfxuuw0Yd6qHBnTzsCcOKaAD7QnA
no0qS5lvz1JYUuZrdMT9SGd1FzlfrbK8OT7c5C/PGcXaVEc/b0dtTHdny0oqEJWP
tgdDlSkaBXhxBgpKKuG1X9XERll1pBNFFMQ1NAfh6CIyj72dIvCCVa8sOGfrcmmY
5pNp+GenOWzPb1wTwSuQygIsj4pcwj425NsEq1rc8P674lHQR0Fm50QQ1gkDmYqs
uVuNhvJ5BzyDCxNz21dQG7baypPbHvtumTTtwLcFpPRHrHXOTF7T8qaclVDXqLQt
zWCuPc4TBg4NVTP0vP13QOnURlFeB37nfTCj0j7uUtylbwVu40FlAMjdbeTaGNJJ
fJM180ho2jO0WHV9hDQ81pr8cOAFZKvYSy6M8yZlRUUkBnpGzIAbxyUMEbuEvXmQ
plUN68obLHCfeDR+iVScXGU2qVsbX5cGidHQc+1WtAUj4gImYq9g/XDnOkW3DG85
JYJs8k5ZbUtDmhu6/uKdH3TUmLy57ahPEy7Kp1f0/t3YkLv8wDOSIT6TUQwiXx8G
coPVZkzMIVQNAjRlGZv8AINYvzg4TUgPOHhTs6rvOuxR3Oqo064KuScX2QS4lbJ8
w9Pjgur5Zc4x+EuU7EYTyN4y8J10lUpTbA73/HPrpBZBr+o8C8khaKrqW763xraA
WjGXKKb8r4ORmgiw6HMpvuiYnEe344wblsRiAM5C6vHeoueIQBl1d4jR4Sy1dBIn
p5P4et5SuRhtMd3GYbRD1oxkNUkFUgQSVZiZLyjrLDQOsnxYB08SGY33SwhPpL/u
l8L8h1XQ3ZCj+gYSDrzgjk7AQHmSUoW9zWALatw99gSuranLT0h3KPK49mLtlJn4
RLH93yDFOfOF8E9q0n4+weiSaSk8A9HrfKjXJJDuulsLZg4DFWRq9y9GA5nB/pKj
gg29uUKXayUcxv7vTeqm0bYAs0jKkeaQAYheUwuF/7AYMYBgIF8bwJA7ivMybXxN
+6JXJxll6ALQ0ff3bqUACjXHqdVn/hQ+/+kC6XqIWbVnOo5GnDhy2OMt7iTjXQVY
+tQw8TIlffwQqRVxJLVx/++wQPHbQY44NRDuZ/4E4la6MoDYLdi9fzd3hRx5cwce
bCpLEQO/hmW5NTGwzql0KFg0JC1/o6hjR2AB3ZA71Gcv2NsWCnIrPNI42WwEHmjY
UwGeJjUlvOL+ykZ+iF9KTkDHOBynEuCF5pRUIne7JHn6xQLbQ6THzDBmLPY97JSu
W4u4dqi/gGjKXQmWBQ2Lo5HiEomj462sEC3Kxdn2nZq/4Oaj24w/Yu0iKU8xXPny
B8eelC8d1Nv7fhNQp5X+wCnf4TgOjAfVURb6p+ORXRp+rQ0aKNckXu+SaKy1+R09
VN1YjLLlx9UjrbCd/jk3oNXq+zhPaDs0XjMCnbFVRS3l79mDB+tkBty76pbUNe8d
ib0tZqfTQFMiJDUN2HjKJ6C2O9phYgdel6iJgkf6CnuSMwTB5lfT9oCch3j0QO4G
AdgpvlUgrI1qK/A8pUSWG0hdal/9bBzIIoD26G6H/fAHRznpkI1IhW6wnJbWlXsC
+BwbUXMomwy4qWyHsyEE3RAcLFxkCh855jpBq7gen9v2qnkYVbX072dCpo/OMV4u
4j5eWCZuGZ4waPYaj1Z2mwZHJHVU/b5xeFUYta48nbLe39VBHjyPSSOFdf3PnpvP
au70LsMuzA4t6y5i/QlYQsfKoA+QUXjhWu2Cq++KaYlKpXvYtnO9JpNkQcowd0Hi
iPpztYnOtNU607H0IiR374s5Id6+0Rna2ZDdLpM93KnrI9th/oSLucPibzUUaWuk
dDPrIbiAJhyRnK7mgvpXhK6jlSVCVtx86uA+AMHPHNI9VslaVZ7CcC9K3xCitapL
GN31Xk2LhWV0UzMK1be+kt7DVPupgANy9DlnfoUkrFHzsZ0PpTOKVL7HEkO27CWd
r2PX/FgkNOmIQM05B0Ip0Zc0A/gYSck0e6hGkw9AcjIzCxvzKUWtVm0yVyHGKv8d
Dsp0Ts9KrTU+G8yaXu8gHGQFLbWeBYF3ZcxsSXrpsL2SE1h7f4PPUW49rYBgszDC
z/K6o1FcK/+TK6ZYJ/1tSfe2OC3eY1TypbR4zGpEUCusPEYdsCMVoE6PDndzp5eX
r7COVdhskUZNWgw5llLSIDrc5peiM6FSdVNzgj1duMM32A1sQN8XRvCOnib0KEz7
y49oAPvgA/F1/AIHgUAES1FXeTdsbbYbD3/XelOnHEnthgbCD79JFlUpWtB9HGFo
rAf9YCuswIyx4n9O6/GOHZfUeRgyJlf2yuCjW5zzbPolcQ1UuuGgfCuhebgy544X
d8JD8Q0ae6RcLXlX912Z3sdy4xlWKRsL+040UUQlHVKRcA2urlbFiTWJekneAttW
JUuFH8Uh0tw8zW4UYQBFiujveV0Xit2cUV1qzbINPLVIekfu8MgZe4YXpbVTsNwi
LUj8K2L7gtFv3sYy5E23mG+od8xgElJ1E2lxwRPmMjIniGk+1AjZBR0P+DOUb8pP
WlcZaAhK9qXm6NDny2eyWv8RRPIhMC2Iu9d1atgcia4s1lVpJ4y2EpGUfOj2sR4h
g4FBIk+SDYGP01dlBKd4X0VOyHxxgNLRV7jC19GFyvCjNB9LBF0hCWUs30DNzlh+
zugII+L7TvkHlVPZhR8cmO4uqaQZ3KGhjPHeWYaQ3KuSlF3PNepNQ+T2eZ6w0mOZ
QMKxx6AsoYsCoZ6eYNA+3xXFJhDwWpxBPG5iJjRUdJCAWPlklGwCbiVpkL+dipGk
eqUQj0TSXBdL2Zj3nWI9vOs1gvYqTjppy2KtKnyKSj9rAAPvSkjTSlzPasjJmIrx
fxVjvEKc0FwnxUxE45t0/mHkomtduFRYlMA43cHqoZe/rU5R0yfQpSxooHrDtaT8
fesGMs20ffCLlTFbrSM6ILqxnIhT21SJfic0GjFeiuVMtcMV99P90ykWrbV/DU96
Jh6wJrv+Xv9n0bbYeZoeBd/7FxOVLbM6orZu+zfJrVht+LaEHqtKpqxnvr2uOWlp
IhelkHuCZuLMrMF3TufTmEk3i3bHwb/iH9Dks+8+XYt1i8/2Eo2pi0jkLRhqr/rh
mQnacKTcrfUYkUj5nUbTZjypMgW/DWj72fqoTbLmGFeBsSneWgWFj556/dyCYXff
EsVRb7SDrGUEkRsyoNSAwd57ctp8VjCfabOwNIlsPCUTlFhoxfpKHI58veCCSHSI
jxRpzsR+3wBU66NkqK+ATDexrCy1E5elthGfxoFsINuI/UkpeJmJhcLPROEXKlGI
inuW22JtSHO3eDvjDK8swwdhbIbLKg847OIQczS4oRV4pm9DyjBvWzIjZkxuxYKs
KclmDGiSraKNbNd643E6JoHtCXR312XYY+sq/cPNpwUsElWY1kjfZNscYAufwtgB
MGXf+h2FTAd1AQehJgdM/z/zgZXYOnuA9TbYTIXNG6HrpoXV/ZtGK7QZgWB3R0f8
josHaIqSD3qAIxr5GPb0lT/9nr5a3DPj6BPQOolgOlDg6TXEcd98/lJ5U0oYI+w9
i2GsWQ1Vp+gxdHPaXYXJXLcFfBMn4tDHtrueSB4n1XTvBaRl08BWc4sb9YVa0+LW
n2SbYbX1ZYXXp9boCGFYvX5gvHwOnCLT+0mYYv8IGaCvVI5IxS5PrzolpZxtQ8xB
FU1BvOP0s+CqmGUzOs1LGoyCizAVAJPQoitQTkITTLyaBILuIQLUn0LCqAMsX7Cl
BOZWpdKMPtNoZvHhHx24NWDE537wyJAz1KZ3Fy1btoNPxLxnKG49+jWf5nEqdSkD
l3q8tMbFgT2EicjAjKsuiOuZRQprCqBtQGllyf53oGyl5jcAq1TRw4O3zuRYyPJA
+FwiG3P9LaauhrJUKRAGO2C5zEMiukNKjUXaS05u50neD1pN9nDhRT8Nzpgsm3Y6
Jca4BqCZNxqnEACVWLIz/fAbSJmquMZaBvPN570iG6NupSGUz9yyxtAwetUo9Nu5
IT1B2MVgxnIXxXsFginmaxua2RjS5d0SWg4KEExkBzYTPS+C4cQuOM/YOjj9LtoE
5gJBOXZCZeEm9LZScCXvwsam05l982SFzJmjHWHqTmGxzyIYl7UtBKqBiv0RGw+Z
PYJOTdg14C8aeLcGps+jQQ9x8zYC+wrlMz6Gy0PP9L9GsNattTMOxGtEpgtk9Lly
eSHhaf7hWEdcon4K6OwW2HqRAI4ixOcUTXGhxdtYro43DwJdpfFrcRQa/M7OmbVA
x+TVDT+CkqCAfTwt7JVw9TDQyma08PS54zJDka9WKiAN/u65u038zQUxM5BE1ZcJ
63UVNkyuoQHeChJ0WleboZR0YRyY6BOJUEdAvECKrXnbTct56BrdVELbtuCkFbWM
kEfgo/KdiRBXTdQya6qt0tfEfwXuiZvqrymgG7HVsOOtSIpt1EF2IFH8FcJhMe2C
dtMLoXYV3o93zfaGPycECDyNQYWDoqKUtLGRPxc1v/Ix2GAia4RYCWlm5B8QJWQ3
owp0inWlGzq9Jezqpu1Wu56vDbvMqA+UpIPpdz5qPrJnkXfGcuuNBIuuhGKPun2j
WVyE9mpPyBhlj9gR+LPSVo34KTz3MlLd0Z++Q/LtRszUyONDQqabYjJOzFWFVIPc
Q5ZfV/fzLks7ch4Ih8al1/At1VS6CxnqsGgANnaxym5Xm9SC9jT8bxGrseuNu8mP
AW6uJpJXXkv11YRI/m6IaDK8kBetliGcGQGE1R5y5beSUXY/4sg1LrKmeytEhK1O
dZBnqDFUAff85a+lRH9MS8Ao6GYs7dgRJYXjrQcOqNX8HL7++k4nZGDUaAoMIbFu
eHA33I3tASMkd9OwTlrtGDlB0Kwe/lZgQK4ssTPxbztSjK3A6Nw/w+z5yHwUNTh3
F6aj5IYD5VsacOPbLWBS8JuA4kbyEpmcrZmpVzVruOOL3pqAfGVzlMtZChewOUZ6
5j1wqENMe1lukGn19HcvrAtsLkR91YNWvnZ3T/ELuxfZG5iyo4kJKy2OC9Bu3s5W
+5ft7Ta8gFyq124c7KQjp321bWyGc+DJ2jBFsd0lpD5JIuqM6DFeJbahBIPdv2nV
+hNvIAiw9jwj1nrte5euROdT+aW3hd0PLJ3Ru8CYn7OIoypEVRudBWDrgmKqZOKB
NoNhkEN0BQGYhX5uhVC++OCx4R96viRWKR5oSKqpEHtZ1lMtv5sUZlsCp+po4WdT
fwlnYtR82PQfm3ngul4BLEp9FPhXK2pPJ6BJczEATR6rFTisr34+hG8ucfZFpvr1
G9F+s7jtRzCSWceZAa5IcaVN+xJUJ5xZ0pLqwnBWZUIUR00WAZL4jJJysVjSBSSe
kS2+mbnqY3ZjlqUVPLRxLtd6NxHC33O7PkvBPFe9cF+trQLXJ5fNoYP99LIesE8J
q3uW45zm00vl2PlS7Q/6kADrQJGZdKRLpRG++WY1qX6KG98M8A2hakj+DpMbXDWU
Xyy9CG6C/w/n5oY2rhCXRqlV4t2euekHyjlB/QgGpzmjQi6KEJVmL75N5CW6E1fx
1bdomxuZL5qNXT977Q9aFhug7lFHPR90SuqW8CQsSfXIjOJWHNxuzMZ6D1LOd0pI
k3AHA3lnC+QUcv1esMO0KIqDncWgPBx9A/lfYlazwjmTRyjkmG4MYCpjpq1GB2lZ
LQFSnEkJsvdjf/YmWQLSpKAXdFjToCRd6igDQsI0P4SDNH5Uyp5luqJ9v1ACUxxd
g8N9YG7EaoGGhkcUei7E+9g/UCaE/+cGTPac9RLc/sEMcQLiGIp4NnK/oFwzIixz
psJ8Vk5q2Ry76GPJC/DKXBUSBuJkb2c+0QJXOz7Kq1GUery/jewqsGqjbeUl3kYJ
mS/BrDs9Z3NVJ2DUOKNziq1uFi9XcCQFSrJRrC7O7hztOFjFOai3Jpkw1jwxkPBw
CsrTbTjfoInNlEdDfPgZNI+OaaVmZVJUfPQfiRw4m69vHTIL7dXuaUVVWa8yYI8Y
OWjBme+GuPyyfBaVVn8xjEtPVNrLaZH9+kteeXS3btebmVt2YeQwybRDsrHcLouu
SbwdisJxNbvrNkMMj370HuC9zTN2J3oIqt8b0G5XmiAKIQGlZ9PZsVsZB9hUnfMw
vRpX2K/lrszIGzvMe1AmQGFSDn0Sk0KGfRikDw/+1X99oAXuowgmJr0cymxGT/N1
3tQa8gNHmE7W4IiMJ0kwloZrA9rq0mbfaokRayRmL91FlbgoU3lJjxEOWPHBFZhK
Q858OcXhml7Oa/BYC7uuQXPn1LAXYMChnfsqrb2lkam658cX12UIS3dTsiHQOORN
JFacixoUOqHE5lQChuFl3tg6QceukyRYz4uPqi/uY+f/HmQxtoXixDuqBx+V3U6p
36ITl1bEmgjusN6ENjrrLa/QFX1KBqwlcr3RGSwLffyO/mLtJuT0a3P6hrPkhXcw
EdPsikcF1owApxRbBNhrzYK/rgDipTlnARjvNlP2EICjUoeY+zUjygrH9q2rZe9I
2UHFM9azTbAy+otfjL7/Ghom4Cy/x8eEK7SBA1+HlVCwtNPok2cPuIzxvWc7eYxD
53zh9KmhmHRM65gtigdxaNGrAybraJkijV20vAi878Jf1lHVziOsiLBN1fut2iE5
kgC+Rk5vUfHitzeve3rEXZV7OQA+ZaG2jLe1JqCawzb0EJ5TTHaHOAmdu6zfCK3D
fi2+SavNxImMnQi8Is94qIDf8GvA4/IRKlptUnebx7wNmmbwltjOGT9DuimeUyLL
OVJ4x4donk35q1C8p+ywgyYEDW3Lv0TIQBYt+3yD49ddMJSRIReN3VQoLMNakSVU
+F0PuD0yPDGy7P46rfx8gzrCDpJzNf0z5xCGofpCDwq1mE+O1TVO+YGvmIJCZnT5
ccsWCyoI8E67WH2yGmNHJcTFQIqmsQ4uDNnbvUGMvM85UZYqM/q5t69HPhJ91CqC
zuMQs1VyOLwmLJl4/XRdSwR8snCjNsbr+jZW4Mm4aesUWNyKcwrx+/6flF2bwbbs
748W0DpJnGShcxGQ8HRS+sg3q37mcVL98wrGOVSA6veXfLF+OY+zrWpNgZBaaSzy
vJFdedQerUHhmS2fbaTGwXmzbGn/MWtCGSnpEwkZMmnTb6d6+EIFlGbNn8U+nPSg
JbX42pr2n9MBY2PLA/wtRnfgNXg9H/O4AWXtUAMrEqqwPF4QRFN3M5K2KrsVT86m
LtN7mCz8xmWA2yMmhNYw22suV3qgprdQLJaOFk9crBxnHqPX0pfK4QsjJ39vZCax
CPwEwKMgyk3NQjCWnnTUIlt4nua0O27kJEIyH8o1KAB75NBjOdtnnS5105r+zU/W
AnTGaptrm4+WjYuKwQX2oLCvs1kJwf6de/caHVvoU1KblC31VfUibbRe33Nr4M7T
Kd1h8rSUAXXPbVNcgb4fY7/d7B8cn8Rqa67LXpKUQISpkMN3pNHh/klv1nhT+lfl
S/sLwzDAgGL7m+rwTU8ZjgwaCySMW5reqJHbp/ZR8UaZ1DC6cB2aqaGQWwS30UKD
E3mpOkyXgsKgAzhFy9KUPpyYV02uGHZ4SAlC9qWKAseLI4T33jvHzneB8HKXjV0Z
9schZow/J81DH3n5X0kzbmoN5lxth0lXRIaSx61elJjv+8JLKqHnsY2HK6TbucDf
/LM2Fx19mXkM716MXz0qjFeBuY0h5JLZ+cT1uDoDiDw/klLUU/FcChyd4FmAiL64
uqnkkK6QSdpevzQyPaqy+8bR3X+JzwdA53iBOmoDRMGn7GPaefiOYaxRFC9ucsIR
5oayUEX+dKsSXJIBxmCPVYJI//V5algpEhL1iy2Bwl2WRKeVPkVFMiMu4OnSWjDR
2JUSMnr+wXloAttBZAR44HooxG4l+kTI67mA3E0UacNO7slKlZthHwOQ7ZC/Maln
udV7jGatO1yt9OtRmRiFn5qEg98C8KImdJ+Im+U/12r46FcQgRsq/ucXx+qarhgq
q8UlTFA/0g1iIwXstLBu3MZuIzTLgbM8EUuUqx++LeBeSCqc+Lr7h2OtVjzaR1fc
VaLBKEv61LZnXfEgTMaALHkk+4qjioIVdNG+fChhBDxevdmyz8PIBBTLEDETtLiJ
XlW2dlxIi4f403hjpyhH+qG8yah+rm0y48mxAbEgrjoafcbwyVAVWdKdpT39DGrk
h4YADJMuDc1xyTFiSLpYP2uWMSpIeLAoGNmFswR41HqvbJzVFnxb3ADkJozgxFEr
wFv5XOHyIcRROG7x6G/dhzkCTox8BF/LPmebCK0EJyrbeaPER8FiQo1zVYcRRwVY
m/Qlg4Qq8VADgyCxHj+8Tk5s95zKjLDCo7VsYODvn9b4j7a+jAC5S+yh5UW0zp9b
zt+hmT8j27k5odnjffOQN3KOzMZCet8G1IWX1NEK8RktqjZrt+dOkngg40Bj8l24
s9V0slZtgJEP8WEjt3L3YBbUxxByChaq0lOwKv3BPCEaIXpvIqoqnHk2LBinbmHA
aIKteN/yKynhh5re7V3+n6fRaIK3bYkvo1cmjD4PGzKjz80mDcUk06H2HI84v2um
acwkmMyaPgSZ5EHWf7qd4ijR4tL4Vgpoxh7QuyqkEMdTlCEIh6NC6EdLefC/M8xB
2zf4iGJS1EuXvIgQxtzSr5YqSOdECQFKUzBjJy0yrjLmrvTA1Ymw4Nkxz3kFHO2a
HsUTGFacy1NUC39B63gJZUOwEYwgfx+0tAMnme0LHDng9B2zKbMJOxN/h0iK4LUD
7oagbN3Vm43qjBfzK1wzssWOCdZWST6+z9kfOxiBL7Dx+T8I2lVHdpBD15l9pqMU
VU+HqtRjrpsFpy5Sx+gPA/avh2F4qdkf3RbF1MYWWPD5nUBK/Fv/0dbqOqzAHYwY
8iRRZO/wVnTyVI9K5lQ1FX6M4k+pbZTV/pdmHVkyWC5DPdriV37YoX89TflHiOvA
vGJHlqGFm7jLQryW5LDR5n6UaH2IGlNzB/PXeo3M1pzBYThgPNQTvxzyjMohkA/f
4w3G3ajGaOr58up28bNwAAlmWAgXcl5P4kWfPy1mUOjGJKxJ9KMxKtVwO5XQHDaJ
3fa50ic7Xgk61+pmzmjIrTJNpnz0SoR6b6xiO6BWW6pelHSXB6XmAhyFU2ZNT3+e
0cLmnvpmfuK2fKsJk43nHj34iLIguqkPGwwKnTirfGTIy/7vj2Lz3HnRGx7oCNDW
zdXRM+oLkVAcMMwWN3LMOwvIK48bbSPYxrDD22ebMls9RE+sDWP06Ct8MkWMU7QU
EZ95/vbf3K1lWvbraFDuTiTSvYLMnvgLC4fRyLtE/xouhAaYBZmS0LMmWnL0LLZp
pThSMNT34rLxJRZlZgnwKm+C83BbAEgJCRt3skXywlrqQFhpKGEGHvww8poHpkFw
+/W1G//S7iku+EuqlND7t7QmlGnzrivBbwGOzOrHtyS4ApiS28PYtPwrQ+7JiP9q
g4ShGVa2k3c0RB7Z5Y6D0LYksN7zs7ddtU0g1UJwqgCQkC96L3TUE7FLUOwtbRDS
BgO43PlTCRV4ydxBkPolqn8D7N4hdyVOCZMJN2kaMz+UqGg78AFWC4nbCFcW1UDP
ufDWvYgeHrInzzeFQuR0S7aNZ4TXtue/gAGOW2PvHAjjJZUq2R+vSkR3p68I2EfK
h7wF7+hsSqecVYWzQsao4dMwETcxRVH/0+N/JK4fQAv4wLukkBvrAwT4Qh4JLfff
8iYC4CO/orNWDhDcTqxPEVVau4cuS9y0Ru+ZWwe41fLhCn8zyf5LZry/kK5nPoAi
QagoMuC6Zx2WxgpoSExozfJG4seh0U9sKlQ0Z2rAFvFsgcZr9QN5xPSbDKLg1HQ+
nLKFYQFMPUEMm1qCNaFZAWEDsuFwx+5kPzxmRrhjhDz+9hoHWqhaAUWyuDP/tQRC
dBi5CIWceMPbI5pRjegNFMSicAJAK8t1i2d6R89KqXuSZJXbY2Cyhy92ZJqFBvXY
yy/2l1JNDFVO3Wwz/c82OWX1GBZ5MYdSSJtVuJzS5xYlGWkQTm3l4vCcW40FxNv9
Ptl5E5uFQT3Qxl/iRm0yd7dD7NWMlJIcwZaxdrPFLkXGY+AGYtS4PkPUJdOkPqEm
wuZofsSh7YNTNJR2HS2MIY0jBjDgH8Gzq/3OBT61pB75HTM85pDObQZ++sKFF/A9
px2aigyfLXQCJuzrgflLW6I/7Bjs5t05/S6jVRjlGVwU1iwkXftGU0335/42AHpj
DvpbPuKgqGXK+BaB6dXN+DlXcmmiBPFdT8hxbTB8CNrVnj9UgXmqqVL21QJCTYB/
X5cMfqb9ZD212j114Vcf/lubjsihIhBf+zWuWc6fd9EGNG2rJl4+rzdy4QND3QE1
LIl/Q+xci/3CoizDpg4IllVkEC2w8U00w0ad/6oNX+/JGFij4VpxtrkZIThK04Mt
GN2/LKBasZcvfAI1j79eCMJI166LLuzro2cSUTibPKqLtRJOsdJ+LpPqV2i44IAy
OWwJappv3tdyOZEJx04qLFoNgOq3cfP75gJ5r16I2UQAhRwGQmgLUIV3ok849pDf
1s0u1+X8KUYXOOfv2iFCOf0l8sDHu7hsp5UEUsYq+ehWKj5c5mk0orCKmkHqsVB0
0GNjaMq8bYNpbafzxxEUG0KMTp51k+yFXiPLMwpCSugK0bDy4bUjDZP3UBjAgvIR
5yDSR/5QjgP8sxtIR7L/1O/49PGLTybOkAO7qPGqj4RxQeh/EqMrEsVA2EInKh0Q
eHI06pheY0QY7mwQ87pPm3wLilmbvA/zakZ6AchQEg8cQwTlgWEgemYNMVnEEs/B
+aRMQEoHHiFnbcLtkzvtE2ei0yn4gt2m4vlR67VF0e2h0njKQJfM8sUKg6iTUSAf
RtVLHw0eoBpdi90GQOEHeCAXt6THXJawkuu/qfNH/5YwQiR36AXjnOcI0l0QiKis
wEPWdB61uO0TMJDnqP8TLjCA6oPnLJXSFbVe+C2mJNQXYt2FXskNMyU3NO7L0ZUH
HwudXdTxBeLP4B/lVqZguhPNPGGruxpPcMDdBKDObWWNqyvSdgVCme2eUZwNuCBb
M1nUojyuPWLT1CwIQvRSTsAM8JtFfqJCtQjpOqZMF6xHqZGu0GoZ4xfvHt1O7aFx
1DQTBcs8LmFThcOlFzWvLHIdFSAT5sOWl1WLQi/96V5/kphrB9Uj83v/JOXXmbTR
3fh6dElaTjmUq5TfSs+oenVha5tLr5phuTwpLZGT3IH3A5GcruvlWPklCuqh5zKQ
09DIFcGkRVcFBtRB+ZEwytnomZkQffiyrUYKl3Ei9YIl7/UIpcPdv7k65SvUARdD
O9X8Lw2JZoE/OB9q73UII8OAHWqFhpyusFamzwgFJk544ta/q2SOXg9oHXxYgX6B
JS39nIQrvtkt6EJvDpWOUvD8jH5HL4vbFr4LMDIEufmevo0DksDRB+RVZ987/kPw
dwPn1Mtp26Ig1Q0tQe77NLrjPVVeeXO3BOvg0C8ZB8N9977GYmKKqMqlZDSy9DEo
EpJZTgFtmsFkRikr44LgWqja2j8ej2TaFVS7/ZFpO3WGkWLzL6sKl4u9I/u786Gh
S5S/t0oB3CeQzlZskCJb2lqrjlpNMO28PLzBRit2acaYCW0NCPDatu4OSLjtuI4n
di0layxwlWfgsm8e+C+YqYqmZtuFAsjnxFjDmyjO4FNcpC/Zom87jEZYm83q8Fti
XC+iBSHWs4Bacu1ZR9l4UAJLfT7j0btpZhZVAqE281VoBvNnV8RvbWDyzSh7qR/Z
TlOaT6hFUgxBZq1Upv0KuG/HhbLBDEOq5i1uzitx3FbGtchnyEXyFYWmYQ64h8Jk
91Rib3C2ygzlS0dvW+dIZOeZvMYr4eK8EZcjqG4eErfbmBYSV7WDhyV76ofmUZU5
BLa4SZ/MKWGtVdeD+gr4lTYVShNqiITb6BbONJSgAWoEgH8B7GFq2H7CaI2UyjZ1
trwgcKDWcLsUuNYJ/6OTCu+CbuKFR+02aHdVfzJmKlkvCzMojY18XeDB5gmLmTNy
8t/Hu1Tzs1brgPPoUdd/wfUCwsOsbUYJ00lNMNgqF3gsu5lzeSfqNMgyiFV1Bng1
jA1Rj4Di3GqiAIyLf1xQIBnSx2ad3V0LIGl1IIemv/kWFFmzObmKHkZqK8U3eiBL
35S5P33R+wq5ybWqZ1h0JyOiirAMQHgqVIObNxS2HMSO9vIp/eKBpjq6yzhWkwhM
j94CaF++tBOxP48Bh0s1lsyXRXMZp7Jkkbt5RlEARkHOoetVe796Z254tZjdw9Z6
7cIvFQSE/BXTE2bigqXmQjW5MFo/UtiyVmY7U1ZKBesBBc3Yt+qy6F5zZc890hWk
/tieAkpdD0YSSLse50jfA4nj/gEqpwEinYjimjb4ey/YRmFiCHQ/B4PIRRqZjH+L
I6iTaNouMJM/XtGRSdhNBIDntSmk9SlA1R/rpDbn6+ZHSE16UWpeMGP50/gSnXfe
LI4LkRcUQjY5tkccHI3e0s6YCTV5XOjo0ZHnVY49SB2r2WYA8zhZF9YN85GuJFQL
Xc0eIgGE8JKpPjLVgvQHSJERSfR45jb4oXT092094s7yJVuUGhOi8+Gby8t/Ixt4
Qt8GxOLXeO03v8AjOGB9kwLvKIak7x9IaEqhbOmdimaonOG80T3Q3Ygd5PML2tGC
qsxffg/cJ95lmUxkgar6yojwEzHTpnkitowa9/6XNY261YbIEwqml0SMKZ9Y4o5b
+7OHajfCzhB1eD0ZPX7c85rUO3OT8AsO2p7wrQeHWU/bCTfeKQ9dbZA3i3aKlGlc
dQD6H24uiXgHYjo6tPTadyYsowbO5Rak1qycDPW2XHwcsFjh9DXGIdh8OJhSb2lR
yZsYQl6FD59pwsrUUyG+Ws50qF2iRkOT1oAUAHnObdgkTbD5xdnUGvvx1nJ4059I
N5cE21a3MnDhjH5NvsxMgjXKy9Nc0Lwk0MYJ7owQaFExHXgYMGdhDmoptR3SJcHk
WhEDti60alfvhuESavnBtqgQzQvlokcxxaUnOCr3tq8e0j31Kh0gKHkMLksOiLHv
W/wlnWoSOuAa/UjSyMf88uXfhItK8bHPD8QJdUzu4u6q+avk0OLb5vqE7OmPiGgP
iZ5IUsIdjk63+avXFT/WLSNIKE5LXjy9e0H2Ua5e5wp51uemBFeSKuWq2RNlymgU
vLCZfxgVeiL5QGQRgwJ9eRog6ir39LQguWqsN2rxNunDN3bd0gF3K/9SLrEFwKEV
AuANOpMAk2lP12JCmAJ5BOXL1sHNGmv8PWBY/I+64EHm8WFRl2EGBwHQKq0UV+mK
Aua0hFfDZXLaR4gWejJWDJZWBKii2Gw+nx6pUUS3pKjqPmFXFgSShOHhO0Buf3zW
rYTcSvPCcYchzGzh/I1Xneba/6odn/XNYhCkCBZr6W5PiPU3zfs3qPgxHleroYA6
CL915iGwktzXugzTbzVtR3exasfGmGTpQW7nz+YL2HkXlYVDuQJ48X4Z4qwAuqKC
sGW57lVeqxmarigjjDiD5k4Y+YKUPQRo6hNTUkgHaXe4rtjOk4Pz3UpU9N+yWD8m
qzY4GwuGHiFBqCthYxPRC0dCeS0/B8ND0u2GTXmtM10ywdUIwuM2wxO755bFT8ia
+48aypoNjYBIoCnvMuD9QXfAf4T5qZJTubCOE+cCfD3rAKqd+hvR0/zK9WUaLRsB
IC0oFeBEguELLusEyQsiKlNfBj6snikizu4Qt8ij/Q7MaTnFIb23wE8SKCGU1NXc
viDSaHko5CZkdDAiov4Fqfr6pXGpk1do2bEx7UDI0TCo72gXCk6lt2huVnmrSx1P
rbkApaQ8zTBLjnhTvRaZ48RqvLi2cjH582KjN+DNmBVdzpTygS9ckLviMTcfQxqF
L71tDWrkW/BhqO0iE0ksbAqX199mmSENAJ5IWOgVfjbpR9MJyuYAMdwjwlb2Bgcq
+7taKWKDWXes+YE2s0pDKR6S/6BaYh3Z2BhF4WVAFytc5+3EpTdh0O6tBP9AWM6W
72ZuKiXDcEwC5qjj5SiqH+kxPueoX1LG3GsQbTow3jvhrqisD9lUclPV5duSaaP2
WCG/iK0y84nLMGenqSNIqdgTdqLl0VeRW1VkCNaIa0f+YhPeDjHh+VjtBjHMd01L
5SBOD5l5yaiLhRT7FTfcfqmlUH4NtI18yA4pOnjGE/1BjXFV3yolLeNcdfV8fCbv
pxyxu3mLRiS0tOUO3ESk7XmwvLq4MnB8FOGvr01EogWG/I0a9P9jYAbW2JV4Zm4h
TYc+EOGyNP7kHY5Hdiqa0epDAnCk1jvxDnO/EDVFAcFCBtSYopFpbSc1LgyCfarQ
phBg84wPzcu7na5RzvOTIxANaGY2KYtIlqcupBP/9Zk6aXIWy8rkCtzy0w2SOz86
LszaWUw0BUGxW91VH8Pp46yqWiDpZ3wsoFPPfZiNiYiZZbKna+uudzeytPGT4pCr
8+WS+jlKjKl2t6EXDPZBE0ez1egozIPx3OCBHw0/OEd09ImHVR/bseXFoJMHUm+N
vRp8DGHPDZTDCO72Ynt/hR+lbBtms7fldsBbEvDmHr69oz/GbSqBxIY72xi6voVZ
/JgvauXoHWcGYJHcJ/mg5QQPsEIYWUCU5Xoqo5yW9jnf/OTCgFaPeCbkp54S0Wl9
MAfoj3bN/6K1jdlM3Dp5omkJq4My/E5pNuTPi1Q5udrasa/hmwmrKJ8HVBHAK9Jz
TfInL7pGvTw9M4icMkRn+myMyNVhzN4m/k6WrdVPoMMG5CYCcCvfv0SdGpjJHHs5
FK82plm878yLpiXFAJ1MNRk9P8XMPtXK7CcBKfM5QbInGgjD304pKnJMBDFg9LrS
HdmIzonSZVa44a0ERamunW66zca90ttXso3ekhh+qiVJYLsIjpOa/naq1ghwn78s
vOepCwOmCeBBk+P173u17U+xbWmEfh1KaITGl5V+ukS6scWmUcF2LPcXQkFmvpC6
9sWidfs11vQx97ZOHbftPY8Bl22xyyQp7f0mLl5OCkhyCotQURaJqPGGo0scbz+o
vvftKO6NwkvRJ5RiBNE4T98OxfvPn4hpL+92aKkAtreWQ3UiJAXsTHXiTCJ59qLK
2b8Co7xiy7TyrFSqrza56M6cNgbwmpHz0EXlByDAFbeJYUNWH1EnZ1/KEPOvCGUf
cGwFoJl4mBGYwHjrelpAZi4DXOtJ+mhOisuhxFEOnuhlsQz1U+6N14/Lcqjt+075
g2i+mQkdDubXU0f2zMTfxoOlspmx5PKrHOdFHDzIC8PM4Qt8QlsWcQm2pWMDiWpe
fv2MqOxUfFEv/ED8VGJyUAoIRYDFTjldByLlnVmIoTUJsb4ulU0nOPnAtnWLrZn9
QQStw7hnUgwjd5BkL9OGJC1qtSBlX5LfLTRfVwltQ1YNfOBt5RTcQ4/Hn22nw4sS
XWTUaiIC08OZ5YMGXv4xxKxf8eCeS/pdeWQHGkRlOa71HJkYHrNEfp5s2fghBdfT
HpW4Y/n3P47bj5Yk3Z6SJEZ7rwIqYMYoIJphYObXsZ3PqufoL7XkNWsKjTOFYxsa
6rgxtROltBoFmmbZIqn/ShrZJjxM2GIyIgGi8j0Ea5Q1BDjhOlGeDjd2z5nYynDI
evOU2bPoDgnq0wFAnQ0DLZp8kYNdF0R0WX/EmkvbmLyBgj+nDcWQTBSAzV+TZ/+X
BOhLmW9bjWa1JDSM3o7EpVy2FYbhE6hwwoAdlri3E6YqomgOsVZ9rC1ME9ujgxFJ
psIyyhCGaaXa5PihGw/ango8bM9FBgJiYytkWOd9i43ZNsQVBSu0SQrmRP45dnRw
VdY8yjXYR3x4NnDNiHvhd8RVku9XgIWldpvfE2TurVIZRlhai8cWePY+z30bd/Qb
LMVYW7BYUywz6KCK+ueaxtOjsFk/JERrBs0kuVA/XwKD0fN6Lv3RQE+Syq2Q7o0i
aEeHTgEl5FdyGAaOsI909JlKxsuz13Qc4Ov7hqwS6DaBRm1aDgtNUYL0OhJbjdqq
ekHQv4UHm6O5L0Q6biPUlwIujVYfo3Neoo187ybgGedhKK69vkjnPi8kyppUiOBD
37xZ1XawVFfyUE1eIfkOfPmSjzVTOSaw+F+r8xW7Qdsku2OAlHPsWmX+f0CptzrJ
EMGtqXTkl54tMH+cTN507XXAcDwLkq2b9/y/0O4kGBpOJI+caMFhe3NrdhW7I6Es
2UwmxbVKrg6BrjKJfQWP0/tsDXkGLycD1108nba6eAeSwAPyNB39FHsFhoHM+620
6DX+PloMQkX7bjuvFOwaKJXDuR/T7TeCj96qJ2GeZwGfhHtfI3ErDNwlv5vNP7BN
/TxL5l2dF5g8p6G2Ih2yk2P1Pdi9/EI+5AvG4tO1Lp/PoSXs2SmLILtMYxbemhD1
C5mFT54YSm5gNp+qZ61ayYm8RfDHZvEcSWsdIt5biTJtLCuPEQ2sAimpyYs+k67K
9M8J9MO2Sq5n699kx+RmN1Yb9+PI1seB9vVD1NUqWR+uQOlJNdnAWdFobEBuvwC6
Q7l0QMdUoCMCa8DsqgGwgim9K+yTWNxty280g3lcv7d0KBFlG9vP2vB+W/XAFNuN
9gKlDCjRjKX3ysGkbi/HFdDoMAqU43qGAATVtssWVhCe9FWVFxCl53/KiEzYorEY
bP8F9lcjIcBd+e4fLT1DsqsCSPhIBKw1O1vhb6mHPT3dTqZVICH8ap7TlRvHKmj5
becM+KCwTiSV6hAzd0kgUypmi5DRsbbTRW4KYWgA/eBtvIFWf/AfumIF/5uFvppV
rXRv5vKcVxo6NDFtcEKeGZKek0eqBiAsCK2K+LoCxD0AgjnyhPO/R51csMcY690A
iKdh7Q6XkEAIl0CvaQObYAbHO/4Mm1WTsXPfhpdeQ6lpcU7VtKRa3RXtugzVEAue
7dsdg+vjtlWDB8wZz+bU/RwuqjXfPIwUI1lPi4DfJY7k0CyzMhK2rey6FT2zKv71
ZaBDz9U4jy5r4bB2iwaDad8uTICSQW7508aOfJgdc2Db85EU7pzwzo43b2rDFSrX
Wp7mxgRUbNkyPi+hGZxxWFAdFSJDK7COb37GzRW+w6w9u+2QgN7JtdRE1RYTgYqf
DDhRJcDIxx1SpFihSOxBittwTWxJEoXmalmFqOSb4G2uJ3GTDYXJlgexW5gJ71DD
dDzJZ1Y1RhJ6VdbO24AKlbZ+5s7p1MeAOBmxyIVZ+E5bugDn7CDd7AxLxYaInkE5
fl5LeEfMwR3drKpB9hkWDgSKTlZXlN8mU1USKKlvw9ETM+pPKqjxEKbRevP19hT2
5Ju8OmxAT2MjwqjeAvCrP/w7HYhjgQSq8gco3ihjoiLJxbLe9XmVBtLIsYlMn3/R
ZEOT3Hs3JSO7c+BFPf+uWFEqbrTNPh/x61wpfqve3LG2VK3bXxcziCieJmq9qavC
LeGNwZSxoPInxkpQB1MSjaToX9nv0GoqJdU6DLQ8A5H6E9zMKbWuWuzcI8a2J9uS
bIu+MBX+bhfkCYAMCf7DLUBU4YwP40poTLUXGwPXCO/Kv3wnnuyJo4zeMigioUUD
e/kaZDO1PChVTvSR/MS476xBlJtbMxHHpe5lGaqLZBlqCFV2cI2CI9qNX5l0J5Yd
yrIV4PSL10RYzx8qFsboL5d54ZT+zco0wfyOWSnezZIXtNmLJbrrrLFr3cTf6W8l
ZmmIYKL+0JJ6jkIpUFX+gb4xaJFkCDNTBcNr77+qMOMzBXZuMYyFibZUkQhD3fdi
vDlgBX8OLuRZOgF0AGzUxKnApd/Jx5i+z4F2u6fYKGSp3pGJMe8Z6qOnvQ+rqIOV
9cnP5AqTkdkb9T3PoEbaTM7v24LYEXz+tcKBT7hIAIBqJSg3EwOOFKojNDFaC2GH
kNxr0Ss/t1/Z45FjAeluDSguIyEO03UaVGNREpFESerIvm7DcYtdpm+poXyonUqZ
aNndvNSB8rqaEGRmt1O4SgY6wcXZXx0ze33mNZ37ivyF2yzMEj63dlvMx6k/EA69
JBoanE7GWPuD6YXJUfJ5GiwPxcUUUbsrfRbJ2AqItipboOCLhXsut95vf9YYzWTV
dpa38U9qywvGhcC51VOFaATuFpvsvhYzhKu1beEAswS2SqsUMURXHVO0y4Ybp2l5
sXXtPzE7q3rCio8lgmwPJ0QNd2xIK/JQQYuUwF2ueRUBzXFlGnsTkV2rbPg0vmaC
6NfrDkKc/0r8yHNgCIzZUl80uW6v3Bxt0JkbeqMhXbO8j6jhU0d40oTvLMic0klM
Cw0OBiuzuufqI4yCZ70GjdW9XB2lkBssyKNnjZtd8m1WL/HUIlJrzeEIxOWGVj+B
ErGUBuPrvxhSbPL+wTpaPlxT+I1w5u7fFZc6mxS4m2TPRyCwL0It1uVp58MCcvA5
2t7WooiGOG1Eb2Dfzciqk/8Lh91D1dpGb+jrz20o5VrRP7fhUJ4rxpz8EWR0G5+z
9aFt03gL4nIPte5jMGHxo5U/VuAihR1SVvm1JGJ01+uUCOsIxIdaPymAVU9HhFH9
snSOvj2g6Ck92YpICkNou6O2jOxyhsXlo01da7/hVGeDsyw4hW0Fj2pwlU4wZfDC
r4m7uqEnzk/lbjtCIfzYiTayYLrHpA2fSF0sHZe+vyn43oTvZLgd2DUbIOb6LSbU
mxk9NP1gBECJaRDKsgD59IyINi2oZ5py4gN6KgugVBJui3P3NI75yWutsLkITo79
FseB/CwFwgMsmc8ZKm1+YcfylBs3Uxc4y5XqczR8NzscPraTIFrhxua87lVGsG9q
LpckMXfGYYuXay5OZauSinDGSG3x5N65KmGgYewtBLOQNMuH+eeWeJveTDIqmH46
WFeZBMSvriFSc93dnDPRgE+Sw0DFQ7CKl3lQkRq53EOdlqwYSdULw5seH3iVbyt+
ooc9hWRM10W//u+qnbCbMyCJcPnvFG+Zr9EpHK4J6Cai3cFWZKm0JKW4zhRZ8pVx
qyIOJPWrGOVFAPqFgdbb2qUtdFh1sCCBwQjhnH56s5Eaxc9yCaq9hpUz9jXUJMsg
vfl9DPdjaybYCWyNXZ67fpqVWJuAW5AlvXKb1OW0Jaitu3lhE2dFxthDFVWOh9ZB
NTOkkaf8PMPB1q8IsfjrFttebioxq4ggbOkUULrPkf1noO27Up/KhxjhS31KQ5wg
LzK5VxkQ6Dq1dXCtp7fWJA5kc7x6qYQEKQo4nfmQRdXm5NcyXUdnNqBU8gGkcK24
ekGWkY8EO1bHDyHCzahKfGMUWrND/y1FcCylyUGR55y15iOJfjRk7640Yvoq6hdi
WaPEsBezXyDtPliDy2kTauAXz1VdBxb79XUtKZitvprrkt279Ue40/3z3VWHCh8w
OJaF9npN5bRW7shNucWS9ZnJt9khPR5NyVIxhX1KjdSnL8VA43411FoYu4s+Ghpt
kQGVzV545ZRvh1ol0asCEHRMuNMstSuNzfXYgVjy03CUNKKZT8dWDNlTF+OZRayL
ar72LjTFPIwU2vHDtsYc2YfnvPxQlkrU/s29Jzt8Asy7TSGu+SnApxEkwMH4cczZ
eVqu2SwCME/+E7QSbjDM0v8+Sj59bdXm1p/Y6GXvI0jRXB2zxp9X2ZGKZb9R9HJW
lSJ0OJT8neOrYA4eHZq2P5PS2ymnmaEHyrgfeolykPHAIVUpiZtnwsrsfQB9KL6D
OdM+guwvqE2YLIEqeJeNoL1n1gCoaxcehD0aWfk64jLu6fFti8sgCoZYzI3437bW
9HQ+9Uo4tbiR28tj9QNE9BqY9VvLxSSnsRTYofuDKSPrELFqkkP3VNd4DZiqMQjj
ouLyZlvummr/INn/JqfhN0fFWCaErIOFQaigVe7lEe7/EEvFjICRmGpJP+8dZOa0
RN2NJolpxwDibly1Z2neCeUDyeoDHjyEUq4CgriJta3/jGAvVRKG3lBuJiVEYB+8
yx/x2WquAMA8bLmuy3juMozpcxOXCe0DonDwwdoxLTS1Q6sv8Jnw66N5hG50z6qj
FAuVq2JhtGdFHY0YvGDXSEcot/KSuGUKihAaLc/1TW0qUKjtkLvdeLbN68mZDL9k
w8MI3D+C7UfW8Dnopzs4Ct5RkhAjsbsF5O3XFWqWCnGDw8N8KLhK/HGb6QeS9XWX
e2ijIcWetc5MfFVmSQsxtYc/wOLzUqHQzSfb77rYkTwROL+R0sYPpxl5zHH6Z3Z+
T9JeCwZGkigG7gqllfDw6W6CCYEHmyBJk3a9jIws29lPv4O/7a7GlIw5ULndAy41
0+sEzrtdnSzd76fNiSL/HVfWxaHNacDHVAWJNoEBqwwXId5BSbnX6HSXovPLZ7ie
UC4y74VLUrtoXMo5Lq5TbPES04I4RRWE98gEFNCs+FFgnJ3m2encaaAFXuJOwmRc
B/rDier+G02YfYwkl3LhYzCAHNwCj5o5v9ncxIs+Et8K67KcKI4Ry9TlmDqQgL6J
oiDoXr3p53XnWXTqcy0zXicXPTl08Uf+6/YqLjr7Nu1FMXiyyYF4DSm/efSs+fjM
uxTVY0n4ytXg2SPUvql5WJ/OChY0DCNfnVMsZuHVnoLfwRhWZTYksQPBF33ruBRt
AFFENoAFSQ0pi698fcTf8JT+vbZftP2ksXPaGTdkXLxq0IE2Jv/LwFTV3zQZkf5S
CHLpfN4ekj/Rs5gC+ZLrOM2DkOEP2QV7CCyshuUpa00VdNHdJDKLxsCpSJyg4Teh
r1o8Ho2m1IeF2QgoIf18kaH+SwCGeoHGWhP4/PA4MvsMN2VUVn/IjPF6N3hG5aZW
wU+XUuvSMT37SZaEAeXg66BF4j71aP8++npQ7sF/lG5x6guFJUEXYU82vM8bJtQ4
GaCHcyF5cGhbSTKaGtR/dY4uvYaPZ8NV7tucqWOEfVPIMzHvmJiLFg+eP4p+8any
jyTJrf/oYMM1Jpe6BLSeqXnnz3ABVBymSkzdC94IN2Oqw8nEXmJSUdbhaGJCL5GV
5H8Q4WrqM/V/NlvqD6/lH0lj0Sqc3KDSB2Iql+ufVAFfBakZfVwZV2RO4ZEkdYmI
yh3V5NKkrJeK9jNtVmpb5CbdFpBZgdwDAA9fMMLP9d6XwVeu2v393kK8U3s0th+V
uxXxPpMrxLRMOCpoNfCjVjQDP5GxG1j3oku3wF3oQHfXV3XfMdynGTeORnUJ1lMg
vQwb/18hyJcOSF/YPf5wsjPVkKhVB56KnkZsoCrEh7QxJhWc9q9i7e30d6oKbtwo
M4F5+WodpgUw34yo50Eu8oF0FnSIW5IT3p6bK/MXwlVQXfzof3r8tGgaRDQ8xE2R
QSa/FlJYkJetdCvHo6692jtSU93tPfM0Pydl/AyRgI3/Y9blf5LOv4loFuL2cwu1
193ZprEIsfcEyxkRAziGEO1YuEPakc1IRylZi665gYwX7OlznlsU13q3whfSNdKL
TazAg1HCHSMuWD+LFzLNPQLI8bdHQJXVxhRnLVDsiT60k/rw/tPEujUte4ktoU4g
JFmaE5/0R4qOJaeTHm5j5QZrbd/mmNJK48bi75lNeE8bcZVguyTzZGRe8aVNCV2r
Il8hzIS3R2OrTNNULMSsIK8ZF1vbr2QAr6a8FRY7KTdqgqIpc3kMUUwPIvUYmuGd
MV3SLzDjQXotozmK54Ik554h6873dJcaD4nX9qYqKE2yHsVTBD0RKWm0+1DXnXcw
9YUP3AETBbPRH+TMpxicMU7w9HX16n/gaxGzDxLbusiuQsCkQkhkiJOXiHWnadZU
SU+zdF7lgBv9vrRiBM11boCo4O17nbXiAhUs79aSx1t7Pe2mpaUIZNnRkTSLJgtd
zdocwp5nbkWoXa3Md53Ca97PyhUj9aPU6RBbGKKHh+axJHj6Lz7luhFkePy21SpL
29uu6MtBqKiwEwtlO40gyfWWyMmmgpI3NmA/xTwHALvY5N2duVcRaYEqg5JZuBT4
h2HJm/Q4trCgkfQiBeOfUYI9Pt8mD1f/O8VKf2sXlBUwL2m6qNPSbMha+O+YdfV7
5uBqoiH+0Cy0599TviBgli7BU9ZRFzDtTAH0PKt1lC7kAM0Ik/m6r/Ke8l6Xhh2c
xzQnBMPC+9a45f3eep3Y6lQc/halQl+g30XJJdkYu9WQU6d6jMcnduMy/4YLkHh2
UPqrbYYlqCcSvd78BtKDM5jJw1H+ZCutAtO517Gv5Xxn5mBlMTL3MtszbNIfHxMH
zHXYIkGOXqpAMGeIHTM/VJkCkBad0FsNCj1eVCwjTVReX8gD1n4uPvqm4hBwaSCO
3b0s1Rsx1QpEjI9dao6fKe9220B413uyN6g+fwxszDtyPgxJ/KFATITksNoi9ea/
hq5TmyB1MECKHBotOo5UdERsTgotPueOhjZzGV3QMOU08GFLamOwroBe84q0BvLh
AO/kZ5W73WgSHqwITcpuoVSskcF/TpbewHnUGZQGrE69XHsyWMLCBNAYIApC3NX4
uUhnfVlPLhBXm4lmEnLekse6seyMv9bKkBzrSinjjJ5/ATLiA8UqygPS+thi9SPy
3C+wMA05Pcx/Z16G1Qt/WJWAl+lFszxLDD1+ds2D+m1R0rVtWszpZAKyWFQLRXbZ
sjz6H++MWou/69bbtOq5eqkd2fCvMTg5iW2jRnM8kdmHV+An5Z1oMcIawN0kp6uI
6e6jbjlQPNch0HzZbiFcgZXKO5dX3EpT0xqZUCatXBo=
`pragma protect end_protected

// Copyright (C) 2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std
// ALTERA_TIMESTAMP:Thu Sep 13 06:32:39 PDT 2018
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
dUvCpk9wLxXpbmFL0PuFYEOiOVxrabuJ1EKIqHWDnTndAbKnvfUS9n5T0p+4AnTc
nk23jtasgg8s/6xAg1Q2mw8/uchRQ2tTOTrZUAWsPLfVIrSqpxT3e61zfhNLKta7
dYaz79LbN+LEFa8qCZNj7K523nHY7pfBkD+9o57FN7E=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 125456)
mdnfv4lyMQwx3tl3C3eML2McJjYQYOiU4AH5TBgc6wzI39aZmzYZSkZVUoLPH2xq
D1S1XVrvWoqG2tnjrzZDppHqHndjvOAhFfTkxAQ93bcy1eAKqWUupXyjIx4J+EA8
jIwOIJ5fP/Q+I8uAQo6bPCdDd9TaL8GVGNanfs6tBsnT5H2LXll1hYRxvgqjxDUt
SE6dheDJg1OZYW31d5KTSi3XfVFPIVVGpnznWYeWJAZVOIDqj/QSlr68XlaMhNjN
X1ABGeYt+P4TptCwv4Aw80EPzTCTApyUxcfQs9Cj+7wuly6X3+t7KhBCCNWYLhwj
tfuTeCFiGK4ief0HPF2reVJyDzb1obyzkV76LFxRlX4K+IOlV4WW9kJiZ1xrs95T
zaexK9skBRTiA0mT0Rb9dk+egNjyHZJrLHo7IEmWFOeGQU8VjfNaRc+kBp9SmhIl
jxXMKD5o0XiFhkLo/eVpZDsodF1vVuXTktRsEf250uDvfOHuXrBAkWjdz3z7GWd7
ilnLBs+lnzLhK6PKzwN1XbrTAOO4GXs+CCQIVJbw34CstDjfJBveQP3jI1TUo+oG
e5BXHIgelYg6ZsWb088VEk2huCbC/h7JSNU2Bi938j4EupbUrqaao7aREJzpPGfG
MuuGXtgfJBC9VuDX3d+RXbQ97mJpW4ANhjYVNDuwoACVbI1w2jEtVzQLy4BawakR
0ipWPFeWlM+fimutsbCux5sR5lLiVgpS1p9xLvyflqOLpQgIq1aaRQMeQ/CtEHN2
eL48tLX13BcCMZqHJbo0DGQSjhDC9UMXqJJUG4AoyIwBknZEJ4gg/ucspQhkipmt
UuxFvtLoLf06SrLX9qMdzPHnE9wicmZW6pNoPvRcwvuAra4sYjzLqjY64mp0MS1H
MTcmaInNF5NXKNNYXnXExW5aPRb2bMIWx7m5wOrAIQRJp3z+w2BIqkqMUyy39As6
8eQfZHF/cjb3XePxuwUqBxJh/iuGfG+U1NnnjgoULeyRh+QEq4cp6zC5NG0N6CLo
3RGvoSaHuWoKL4jAI348rTq1F8C9Et6KNqG0c3fx6DPnuSWMLhsdBv7XBuIUenpq
siitX/R3BNe2Cy2otrmtg2IGxTcFtX0JEeDIY9/vrRMlGAfjLy+oNM3nAbbAQiDR
zn0hoiXxab1M/hTyDvYIcAmnnqYzkJTIYRn5p0uJwhuM6WgCBAGRFz9t+tVUr4fX
uJCggSu/Qk4jsn7QU7JQpYjJj706aVDy809Fy323mKqIfEBtQwJidMerG+t4FpsS
ktS/4JN5sNiP/+n7/uV3bpPhV8RNF6faHmDHvulLl9f7h3tAXKyKhiTQsUQ3RYn+
PpB2Fnjlj7e6Spl2gDeIOr1j64SXYTaYRlDCmmJmuAY+YF5/zT18PpTarchKkD4n
03hYTWvgFEfZ6AGukph2I4zffeF3963a0c7BVfvJ3rQrMw6ud9DlDPmKcJqr2abJ
qU2Go4uIg0CWdf5rX3ylpk8OBISsfvWw9DUfqhdWt1qiSb2zIo1DpdxjAndfWNoC
j3Ct+TP0WUaVOQBCLBJaC1c+n7MeV8u7wJj6zDAq2IhHVPx7RHwEsoDr2aotNAmA
ScL25w9B5jrMGbCgeb9lRWwic/aTrTlrm5pdmwXetIYxc81yWPagmdGKEtlAhTWC
0iyWf4hiEBudbh+hkuEg+zENQGAbVPI9/iCxoDLxkN29eWPllyvDAhv1yL44apyw
KtEsyUTIObpPVDwuoBiJQmAteLGVcWS/kW1nRRRDoSzmsa6u1laltiisqZxzLkTQ
vqZp+DjDRzY5AkdUGWXwyFymZYPKlKI4cSxzFZqBCX6C4EwNvzqOooXeqOFlqT+Y
LliMqhd68LSSiAyITfTACPG4U/wwmThwfGl+uIEoZhMRr7JnzkaNMz++Q5ony95l
+CQQBrxeqWOpM37FCGJaP7MMelpMbyKhewnWKDAjIFvrfcuWtcquKOqzKQciFu/f
dV34Uj3IWQHRmWzLVzmuOX75NKClhEfAOWIpfntjAmM4lvdumYbkiO3iU/f2sG8I
xuDHvkfj3cimX3uuFEeIwhiXHpz5ZL/eOYM/ftzbsrqflQpJFjMafAmrjrEmLv1B
dqz4GtgcVM5BgSbcz4+x/LhdH8/qUarsswlpnPrPE1TsmGPwDBRSrIw1cKHJd+az
R6UuWiGwOrpOcP0wUWvPQAPwdliuJaXQEaq9Qe2ENKKrAx9m0Ie3f/p8yFmBle2f
BoxmvxA2y1fW8Cr0/9mWP2kzLMdRmwgsHqw4j1UrdTe3vn/p3HK6R8qrssvACLhi
9ms0bz70vLjpb+McYLFfXJQTxbp+p5F2z83UsJ2QgFomr0tIBK3gnIfrVyfaGHvI
0MkhLnNNGIysteSkUE8VSqRe4XzHxeWUHlUYWGR0Iu6CQdRNHr1oy81YA6uE4Hr3
I9C+864KyPFyJ6ktNTGumd1gXWZJ8drNm5xCoQ9QjH0GfsTQN8sjWi9l/pp7fCN5
ZTCWybF4SSEpRqnDosO/yHIPKNGZg5ujyMyO6v36rpd6TK6aMjCpFvVkWw5BErPy
teiZjc0yPpDZOTvGObSBcfeVnM8yz1lZvilpLgQr5pe1+xNtHXXylqgjtqsOWKyR
oUrAU9TmG1nzXuRKUftTfpCuyLeHB94mjhN9vYccsUGVcN7QkOCblYGsek2cB4wj
MGfG0HLLjL+3gSLmt0uz4lFA9hJkb2qAwPQPlRcf1DLRb3O351TV78qkGWcuCptI
/8gSY+rMwotfwbpnvod56EyXaWPs187U368oJufxI8D4L1ZkJkZAQmiHo6XoLBd+
MZVqO9ZnB/xq8JRJ+qPIFrYpbWBI66ybNkysJsTJ5UZOstFv9oRKeRGawY6ZlX2L
yRZW9kmVeAAMtIpJ7vcaz8gzuaP2w5XLDwS8PpTLlx7dOFmy31ayumnSIa/3eX71
+pJTy6Nsdk2E+MTPzKk1vuaoZGg3nyt4cpUmtIBnsZDzM+QJS5b7gwHALDFawbuN
qyKKzyraqrUD0lYBr+zdT/Q3hCcQxRhbFNuUZVWeSXZnaA2mSPLGNd3dmALldHXl
4yfom3/XtIKSjHeVUC88UuezcM+756tLsE+RNU0yTPKZS4lFS4LEEzwODEr39Rmn
R4qA4cGHXDQrkCPxDyXHslpwGlJG4MGo7RUKSWXDKNNOGfFVYhk2KOvTW4WueQE8
Qh1lC8cu5WXoa72mZ/30RUs9UVlQiA0RPfvtFQxHFJS7YU5NnkVHUQ42NPb53igQ
67FEIS8Qf90URXtmpjXe70wnHUxzBX0G1rNqa88P8UPDwPjhuhSmEMrqczyk7Tt4
JqW0yAL6/GGTcu1RJ6ufKIEgoofG+/UC+6rmWZa5ons2tZ4v0iyELYE9yRzRDYKG
bYljsQfPLs1NDHyerf5JMIOyzCv2K/LLKieWK41luQxoDdHnMPGbVhfV0PGZnhzk
b4GVAGnzOe+bgtR4EcYT4eBR+ARKCqP1+c3wS2Epkp53iwdWQIC60JfSX9G2+1GK
loatx/I8oR0NxcObxe2I1z02ct+xm0kwj8CH4kLSMdyHSpbVPzk6FN/qxvwVWh9F
iN/+i7mZeho0G8SsLdvMFVCmHya6NVqKjXCcVqfObueAoQXoAIwO3ghmQODAU7QN
9hbc4J38OXEz8oS1ijB0Yti6jimPTf5ie1BKVjp5ha6EKTaDVtEjbthcnNKBezBQ
K3qdaWys+TYbAMasaAKfpltpepz2xK9P1FbZjnRluIjGfilXAwpkdOCT+NuffY3o
Jw4ke3n2GtOM1j6Shf8M9u6wJK1apA/f6el+KcJ6dnCtjUjNlnm2JzgfGHct0ZyR
xsOAXAg9Lff5zk2fEM3+uJOnp2PH/ovPZ/bW4AnHmECAPHZsxlbn5HNedWIbQXvC
bApwoyAOGFkBNG/5BUAdQSyXlrDYpBIaoDAqPIPNGxB0aWC6I6yfVKchWmCaP3m2
6XBpF28VcNPgwhHv7UcP/vltAmA38SO24tnHixdrICnnDmKUAmY+yGgImHGIvvuz
zQp5BCsc7+iPZ3hcv5Ngcr9ohNJZ5/9UoNLUcMudYxamjQVszPaqnH8aljKWrIGJ
llIwdNc3wWwGuQpWiig8I4QgH7dwG6ylproRxtdYo4sViCHT0UraRPYdTsGBMIsC
fvRPvuasiRNlVzcdR0sfX03Px63Y0Llw9QWukPwmlKBMgQpVSxMUqx2aEsMUDb4j
a8d6p9cEzoo5MnWz9BRbN9OK9NtnCmdlkCqk8VL5a21FDHlHpZhzfD+t3u7WfwXB
dcPJrBayxMJHnwGNiDRAFcBDK2RxagbNiJwFURaOeh5U1IPI5nwCTgvCnrCPB24E
whxmT+ZXfpX7iyfP1SxWevgWCYpFUA1de4qJGqzoTccrNcvKQRhm2OVrQFVR+kXY
WkDOqK/P0MtKhvr7Ka1zo9gH1kdPMpG5hWguem+FcqiYWMpYCx0ZdeoOadJ4hDIC
KDrbpZiPkrHWPV5cDOEhZNLwjwraH/2XxssXe2PEcAVcJSI1x0Bs0XwwCYv0puob
PpycVRvks4Ubn6enngzPi/1VEtVJOoboKNURPAMDzgnrVi3prBmw86NcvQaffkPr
XnC4gPL7QjLIR6BMDjw5SZl/Z0IFA0dUM2jgnJ5hFfBSL2teiyrkaRTiDl2mwd81
0RDzlR5DyNXXjhSR/xp9Zi+a2QzL27G8UBJdCwsHJQ9O1J/spwe4R5KpWZHTdvJ+
JV/FKf+De5m3/7dkgu05q/0F39GsyqDGAb3lGE2nMOvqcy20VmSYFaDEaIbp81eA
sR8xQlAA1rp/s4t8lkVmfV2+FwGnOpyHhBSD13rG+AGfvQvBUw6gw200y2h7cz2/
JgPTHmqzDTQr/vFxoHZ7STpKGqZgau9t9bOFVoWrzdq0Bu12dOTw139sJ+/Y5sX7
GV74LnF86M1Ybim5KVmeyyq47HkY8y0J3OktOsXmgEHHpUxpvQ36GRnhiLyTqhW7
iIrKssPT/yJdT2j+n0STpEsMuW9+WhTLgkDKihpoFrF0ySDfFs+ctBNYPw9nE5tY
HBTpT00wSmX5PqHWrBwGLUNEUkbjVsyMskLn/e9dSRirCQbrE+CMh1pYtHGa10rG
buIBAHAS42GkCqQnm1eBCPZ5bMsG4Mk4J3G+qgoJ06bRl3Awxv5zqn269cizld4i
0N84PkV8jpc+9OzuQj82fe/vMjK9cOlFNbpQWyIwy1OjJ4yC6bmdqQ//ZXKYT1a2
4RwqAPYdUpcn0Bm9rmSwAiCfayFM8Y5RwezWD+MosU3EPPzwRAkoyQ5VGxFrTfY1
infHgjjsQJcvw3mERxqw2JInf3cqlG4FGV2LibzjufaxwiodhztLKEVHkcwoDTy2
0HEuqwGUtr11oIYI9JKjfA0a++tIKaTQk1aMS3trgWQRobHVS+kVIr/Gvd+D5oIk
WCLmnEch0y0T2ma9/L17qznV0u2Q153pFnqABNa0nL1+xd7K5QU43KBcA93/caN5
HzPHOBNOHJr2imZXR50/Mm90UNkuLg9G5Tvt0CsWBVimo6wUyN1CvEcKYXo2AjpQ
c6qwBi4jBEtK/NsVGQOofC+ueikYGLP/SeSpDI3ym+u0MhbJeiPORlZ9qqgJNHGj
LXyB49nbiJIIz0GGxjm6PiZtsQU+lQuW9TMXnPwTlOIvQxnEsMbrhRFt6wCPmH3o
TyrgEsZXf90txpH2CA2uw71eOkIhtl72fXaxzWBQrdeWFsKcO44xi8xW1W6HU3ej
nuImknXjCy3FfrcNbd09j7xVYPokn87NwvmzFVEVKPqNvhv28Nq0u0wjE0qVymxN
VGKZ27Xg3LzBGF+i1VMNXIDY5EfCgKNQ/VV5wsELBheIlbOE/Qyy4isNolxdB2nJ
BA0CsHILTmZEyi17339oxVQY7aLmj237ENVHEs+EkqA+dPS6DWUUze22IIoFMg7K
j/79as4QrYOGFWp5SCwKsNP45/lhrAd+lRYjvHyTHDshSuOpFfiyrHx9e5W09Cq8
O0xBRyU3HyVlMfyEBcvmTV74GWO/pBqb/8LvpWwvW4rjFLl3P8G65IX0UPGmZQO4
mhhwEMhEIinYSm3yicHZNp/PTumOegmsEWAJOqhePPAJKltgNlhDPKekKf8fFze8
CptOAjf/ZJ5GZ8dljnUS+/Ew6BaNXiiRD7z0w+4ljPcaBSPxCc1VeZPYQ/icozHt
0E2G4AlYKeKYVBpqkmVYogC7XDyNvaUoZg+c0Zyf9CUyit7i86WPKDqpVZsKS5Eq
RHQpDubBdqWy32n/bO2r16lpBMX7TekQUQmztTZkHi+aGFsq4WasezxQOLeyZAOm
3aOVyltIVaHeOfPK+bGSso7YTYCHjVbitXKqodAgWjeFRqQfIk8nzqasYvG3V+r3
SXvD+j5l3OP+8JrM6y/KyOUDwXT6vu82l8Pjduv1ibc86FKiXfTkRhYYmAL4uVcl
q0Ggdk+PAEL5bCXMUgto1Y42Z9XQR4ezUwL4pj43KgqjZQT9h8JsUZTt4TOkOcPH
mxeH0jQH8STie+z/mDTDd5PHTPCbLEtF24n45Ul/MRuW+As0yXlNGqgK78chlZxh
/LPocdHL1YEoABRM9AjTiyO4O4B+dsVy/1TSkK36CVFShL4hRTZ/AgVGTVeow9Mm
hHfPbF/ZJpTPCghrLRG8QwoA7ZiKJZHXTzHOil2GU9ESEcw2q4BwhvZKov9wZRRJ
mWtWqTxPD0YTznk5WyMwPYU3gzXdivsqyWaobxL2rl2gYNlkg9M4qAYoGWC7H9t6
InOJYL8ziVq4zl9KzP1K2/rGjljHjb6WqKGDFZufBXF0bddcyKUpKwxRfr/8J3bW
8bJ+zLbXYHIXYRB/5eKP4b/TUF9G4Ym1DMyNCMYHe5PMpp2i9Axs8C1CxXRJFHg1
g3tq/T3NZFRQtvt2CpfSZwxO6TZ9Oj60nizSur4Q7ntommCscGK9c8C59e81QDu5
4urHoW1kkHmW7DHQLvFVlB+6xvW4U9mkl2A/88qDNEj4ZAMjHnHY8XMp+4L9bzfQ
8CLUl4BV2hnBM7dg6AzbuuXbQ2tUC5uU3h6AF3iys0WEF8RGmddPgpG22iN8koUG
WRrd4O28mrII6+p9BcarE/pqeJDjeltKRpiXNSnW1aoSFKFEIM292ltqfr0dFWb2
pfxziIA85JpgzajfQ/BLVFV+Ij1NRj7M/pVNEJAIPxzKaLBxi5+xjl0hRO4/Haqb
2xap3LVlaBM+ExHAtZh89INjhTaLEtlp+0Ik0h0pFNlsCLQ5s+WjSMDu8dd4Q9xO
Zra+R0WuUwkHsnXNoj2mUacDFe6TusyOvxYUEIzI66DDT+p0A7sL21NC8juGmQC3
IEr/PBxIQm6/ry2VDayJU86uFl0O3CbJDZYZq8uh9r72nAdptbqggYgXMH9X1poR
h+rtN1lr2mBW1Db4IqLBtzKh7Lyof8Wvrbb0x63TCzH9mxzsB44Be3cdDnwptL31
AUP2TnUzpsa7NmR+d8w99L3AV0SFVDImdq6zOYzG8EhF9STdK5B3X61Vk8odywhF
CQNaP3ZQ1SfqjF7B1YMosImwic8UK3pFgPJ+MnmYttvpMenuNg6sOaOU6DTZKnts
I+71K8PN7zxJ8WpM90ybA/4jdig5gBTzFxZe/iznDI1u47/N+AdjgqXWIDv5ZD84
C6TIGiknrL3qER8BPdwDuTmoAFVbhlj5fet83zNPN20O0+Kjb0RjC8HkFB+DLc63
TdS+VxQb6mi5E1sQRSpPy+/6bfdgkX4MMgTZ/TpmHyvawJ76obW96pHP9gqUOUp8
0VmE+/jxjKn6LQtg5N+8UMisY2tp7sX9Ur/ixXukf/+dmXzTq786zXTS4dCuxpYr
a2/NKaCJyQ31RoZF0LM9IOdS3dfyy9s9mV/qFKCiGHUexyS+4KnfWUIdQ2RwIO2r
7Q91MV6RDhLkKp4j9PvNK3sZ9CJTLTRfnzCaF2ycu0nbwlABxg3E/GreqrCoGpXN
sos5hiH2Z7xP36OT50NgH9RwTamh84tSszhsI+cRBCmCW+kFKx7mr/Mthr9Qr/87
ZULTCWmWGmuI0eXMre/yw+K11pMvwh3/1KWZ+TJIOmSvz+ElSN5uJEXf4kErXAca
89kklRI83lK5ZQ/CRCUDJ9Om3OJc1USuPEBTDVmWXDWVNkVE4zjparI9Qb8ZTQc+
v6jGIzV7CI2Ee4ajQksEVIBvUvesNIf2qowD2gltKH3xXYmmjmgS3kz2xhxgvhW1
i2HBevFQ7STvsOfh0Rwuwb7lajJeD6Dvko/O4DbRrLYgT0utKWMC+zSE9I19PzSi
drssG6BwEngOUO5iXmYuDaFHBfhaoshlctA3VI/ubwQHpcyqseu51tEuRLd+LUSD
ph6R3y3M4Y/aX54OUxvMlGNJJK4kSzAmpV5ijVbU+1t5AgkEGzmmeYWZ/h7n5sI+
L/Prodz10xA3BcmXVHAnGzsYzEbJqXsR0hDYO22xSWsw/9VU69QgRXGmMSmtrlj4
eRhgU9rTPymIxoCvYNoIWwg5FJXS9oB+o1X/IQPIumY1H8uCOgQQqHcO1OOHkINM
8wDCmYjaAcySM8qL0BIQUKDLCILfzaUQPbfQkB6JecLDtQVUIcGy9wWrCisd1Gfc
gUN9w4GnE+P1P8yWSM7PyssULeLsWMXVUSoJRZYJXvEvCO7R5tF/xHWv81501lmR
mdiVAMQPNUZeQVOOLpcQKUDSenj1l4CIZm6ocX08iqDgQ7x++fEEqZjd99GHY7JQ
78St7wQ6MswAv4rO/wLEl4jQ+H3SN5F43gjbFEwAo+luP2PxzaH36nGNuk0j39YC
PLzfrOz424bYCwSnf73rnbA/++xmoki7ahZ0b0Rk85pkbEDolUxe630XeTRpdG1v
ev0jnpPSK2D8nBt2/H+4sZe0qUaw5P24l63CvQscXxgJvKJVJxdTtmYAVFHvQ7+4
QIYJev61UyBB5UEcUJ/qYNPflxBKCnyzyuWaeiVajMrJrE/1XbS7eFcanRbOylAz
xF9MUP2b5Vfxe/Le2qqStGgVZNDwv9RoMq7FRaqn4cao+Cfrvh8KylFAaj3Skxgh
Xw8i61UoE6HQu2FuHDsfm8/IeKm8UWcHA63yvsacbT8pdBN1N6htb/d2fUWwGqAa
V9BV5htazHplO8TCdF982+WvW8jGJuBGdFR4uxDSwKmHOQQb1/S/KkW2gPfVgCf/
QqhslB5cAoF0umg6yND9jNd0Z+MoVpLIajhFKgIx6d2dk/SrhCWqY4riskboVToV
5o6rsxm6/NDZHdyWpwvkCpL7LoAIdF/OE4cjjFoFT85Blot8TOQCYfJwF/Xl6AjC
vc/TXYnl7RTakoJiwZY+IVH6MNGUzwcPUhQJVHUFB6TRA2vwY6I6T9+QO59hvBnM
7lweLbuGrvtsR2R2mWJ5uE6xr0U3mnnLY9YZd630NIem8Xo9IjG5+PbJ08Motx6N
RYGo8voR10466kUONotYbneKZR11bz8BG18RgPEzSkKjrBzlnp1Fx2k8OhWlmH5x
pB/XkbnwyJQOEXciYlLU5awqxpAGXjEzpusxCxKlfAG0dmzH4TpyQSG7I5rddJql
apT/sGLs9qA96ye6260lmgri/+xSrmXxLeolqPO9Olg+w8KL6rvT7vF/qXLj4wyO
hh33iO2hyge/4MQzfv12n824KGT4g9SiyDqUIkoSZiWGAQ2t51CSc16oOAUSYhG3
J8Og/DcUWjPV4kA9r0nuGXk7lQrsYBBzQM4QP2Ppmz9SQLQ2ezZ0qT9O/qEY9VFn
DgWBTprfLzkNVMHYWNx8J3OnCJ0tLaXjYqujh0jM4wcIImn9Bf8mq1S0hvM7vUGs
PCzQ/65XG1p9U9Crbyxy9t8cdayFjSYD/1L5KVQSc7Gk+3axR8LybG31ejZE0pH3
BpFKzrQvQHXk/kswANwC/QHFjGzXhn4OGOu5C5RmluURHn4PY6VwJjcAuuI9EZia
Y6wcosyh6gABwp8EtJ8+DKgCYFzHzhd0UoH85A73PR7f35hhVoaFWIuCXNsbLpAZ
sCcgWHDtskh/8zBy6z8ZrIK5XJzH85ISan0v8Ppbngre6/8aNY2JT84TZMnmqnKC
XDFnKB2qQlihd1JE52u9+WmeCAJW6NioVAYYnAwwGw8hLBgOcNLXr0tDetm2WQCE
ULHD8agogEsBorh79mGNf+tAv/AIA3Y9vHSe0Qh3IC78bYUYsnLv/l4/wVpGp+s/
ztMsyV/us8eVbROmyG/cL3Cd23yEg8WUld/Q7YQAT8Yv8f+pvONMI9sxorS3IwY7
3unxDaKaImyaJJ+RGJZRBulV3eOSv0I9+suMYfqrkrlQAy6+DdeKZfiLHmVHuB3t
UF2A2YMjADY4R5mIVwbpEUKAoQtRxpY1cfD8n3eJtGhUAeoIoYlmr26IsGp+sMo4
sDfMlsfRcJ0oZmBRKfMrsAyAKigKRw57NEhTTADd3PPAleHfdhGuFQTuLa2s/HUT
Fj7ub2GerSu/ONwkeR4oYUYzb8Xe353qgs1Zh5oDKpk8BdcjLUyDLplM5rnBAAU7
ehyzW4rwpYRBcjhHJubxepmXRzdmY7r38oBmzum+H83tVK7IPB0OXJJpYXZAT3kp
PBXQpc5WeRQ2+O5Yq9bpLKQgiuEsSMV5UV7cZcaUeouK1agdhey9RBlA1WgDyNKD
iB2ScrvkFHHC/M+SOIJ+vy0VGtqf0/voc5HSPkoCf/V+pC41WM3vJsrTuvAQIo/w
h6CHikNrFOJYkqs92QxMaAFYmdpmpAwWoKHzgVf6gNNaKmiw/zrMBfgWPrf1zQno
xOsZIR5eg8GjcyeoN8f8hr2DUZzkVgzzvCe2LBrGY7JdWOiEEy0Z2YA6/CW7WZRw
sJoI+vedVRVDSmpGbjz4oMSLUZK13K0+OJp04JxLWK7jnbwbduyrKeisgYpw5vQB
ysXYMXeZOykWpPJ4S2krLv4KnjwkBr4RZPW/XSVqbZnoOzBnGB3ycNIuiy4y0Chh
o+A54iwvagcBkI9zlPwThrJHpa+kvych/ZG6LSK0yZ6uRCCzqwyz4v7pcYfQ8iwQ
jjbCn2fzs+RludwyVxA8ciAP0K+N41GbYNAkRJYrxDf+6gQKvySIo6XdUU8Nw70/
c0KwXhwlQgV284EkxpotncdZMKr2auYaBDAeZIUwHYsoORQ70i5EKNUGzzgZ2Pz7
cmeMH8j53p7jdMrrzmqDURHXEPpZ2+UFluiKyQlGG2zdd/r7pYaG39BQunKvFthh
FYHtezzZIb9UNSG0Nz0LpPQTuU3XdPfR5JYWg7bpX4gt5t/LcoKVgAI6ri+OHir8
JsdQmxmjPduWhYIQTJvIhZqrEwH1P0Z8sKF5wpl1ifD7y0AAkxlCZGfy1ocoM6bp
TUbgMjnYhGUJCESB1pj32DCPSnFn/MFRrgeXOfu7I3FDFf1gWU2hM0V14BzDV0Ff
HjJwkSPqmw6ANXrWzl9X/bx8KDr+WgOCqdL5U/Y6djvvRvk4nkkOhpmMduPm7pkm
co6sQWJdSOQkPFfV6diP6DzXFiPKYwYYlHYEYrzkIOU1ORTkqv5taeZ7v9jrhSpn
QKn1gL7rdLAglrZCP9trwGyVGH2+9ldfXwL9sJrGR9JYKtf/uAYZF0eQIHxiRGi0
5ZHaH8BdWycNk+KUVRaGdUP7lgsfKiVaynSYX6N76p/TwOxTsV+PT78TVdtIYs8Y
GDA5vMrmOqsS8KwHfMvIezKQfwEw8WL/W8SiUzbaJ6YXq1s/y4rNOqhYwda9IdyQ
cF/mwgucsN6LxZXkGeyvaiBw/9nket5A6CHRbb9EZa5aFI8sTGawuow0NillPksD
RpEjgugDgN7n6y5XhO+QmSoGiagmealJ7+xNAv8CwKVdQxOggJVkrMn7G3R7AnL/
dQSq261JWxs8qaDQ92OuQ0rezCQGso2Jyhosu1kFoChv4cgw5dyDRDntAc2p8hha
5aWzNirfSrvgZv9WXIkYat+abpY/qv0BQaGVquK079macWFaENyYLy0r4K8dTKGz
UABQiA4c+dmI2Ur9966doKR/LiEHorDZZOFBlLvkpCvL9SsKVaAfhXq1mIWHaiA/
mkxWG3l+xiB6KWhHOhbxCi0vF1BYFRKBs9ix5kKrLM+US0x0Kd61UJc2GoiE3Ee4
ZU5dAwWzWzb5oKu2Bh3X04leo5342kE+Qy020aqGrXqNSSQYY3xN5W/1mDR6ur9/
/bOVhvdRWFw8ljNrqSjwh5XgesUNNO5jzV+MuEeXhDS/VXjSh9czwC8aMIZFKCjd
/EQFtYRq1FhkdxBjZf4nwFnlct96wy47WAOwRvEOMklBHXcIl80HurDOerdLjm8j
2+vSuw6ijKPAMpdm4P0EQVcKhPXYhaXcIPj9s1qFk7H5DTF2Z7Lr4B9X5aiMyieo
IHZZWBDkKIcWeFDHvFee+BWd3z6tdTKlrfO8lKtMcb+E1p8eQ36lQKCF3vCRublK
G/MavjSE8gu6BKmVLIGbsTl02czvrbO38Tgn7jredo7mEHlyzDOrHbhySZWIAoH3
VaE0Kk953oDapUSPqzLMwb075ef5y86odQojRW0Nz+g2mfCipblPgy5ncmj3TSZW
S1LJ+3kYOeQ1rAk+X2xt62ZzpOwFzbzbpQPytREM1OO0lE3hP3j+Q5LpZwL2SSOo
VtzgqGyfK/PUX/Xg4pCK7rdquIEdGmRz6CvS8+xcXHbrr14boJFLVaUJDHmyEB/N
YHyKGflGqOo3+8QPwsFTHyCZb8pyjTlBF2iFCW/9r7dgOZ0rHknOzRjyZ7hp2hXS
vASjNRLkLg59nZfdgjZzzgyltVHIYNYm7+WP+WXIf2r4215TU1V8RH09JOAW1qA4
kjcXAICHrDGmoXt9WFLLYGizcedTDeCeYsqEcbAOBxT78o53zkyPIdvbFNYOqjjt
d9rcDPMXQL+XzCB07lTstXyEJhq+QpuacdDvfODvycaOzEpi5gJD3kIrLemuY0kk
ocJ514FYNRElhvU5jRTxM5KQS5jEHowMvF0vgf/t8OiW26B9ww+6FRV05otFiieT
31qc0VAgHnQ77+8wyVNZ44zD3K5qWKB8EoN5OoIZsmIL6lbG6VBW7c2i4jv7ffm7
0yqGbVTUXEv5KNU0C0/vAp8CUUG//Okz6IINp/2N8CzwxOpf6MCbKuY3uyyfNcY3
kmyrNeSHdx/ArVBYX/7QhNaRvyV1rcFlbQUXXOS78yhtvvs4x0BQl2ndYmlvmHd+
qNsIhrUeDBiQzJ8hRXZ1FlV5AVWIz0ulmNvwph1fRKcJv6hgTl58yJK8Uq+azNwv
LXg0EAlHACKfkCl2yf3Xzt1k9tcuHp8Nfe+0zVkgYqlGxJzMLj9tf0lb8jmJ+6gN
n7CbAtPw8NLaKHNHUptul/KWaju2uM9SJhspIVBbtn/gh9pEynBoDFnyTOUECmvs
583sFk9OcsYit74GcliX2Ecnqx/TxO5ZiYMIwKIK1LFLuA+eBgdP2RXRbRwh4Xb5
V6XXXWhL+V8BogLdwq8yhdxAlQqNAkrRIQs1BCMXfjacSKPHWqMhUJDXMUbw8Ahu
QuW9iFFLH2YESfOsqVTkjQryqtrzBds4E3kvzHAICV41MjQd2vs51pjlswmZvYck
EmYE32jkUzvsm8rlSn/D41udWXG1QZzBJWD27heD12IYNeXLasY1NZQ5Nshz72Th
N+PXSQ2O7FNfxDrJfXm3fSx7zel+9jwF9FetJNkOmaCs31l7OYQpoLsgf3Ekhs1l
mPXkcXzrkp4fSDjbefChWMD7q3WPTICMSkwBj2BED2WuYDPxpcvTPwkERpdpBiK1
D5xvdIl3jYVfpV+A/fbpYZZjM4p3LeHV3vzEMy6HcNl5ahXoalTPEHwVYvfJLXqt
z8xN2FXx3vyd0WF23Ys4ZIyj9lLAh6jvqxzcuZtAVKJ2S+coEEOV3oGOsdUMzFuj
i5R25wRrYMSRUMEeEcC0h/DhgQRLR+C2409SscKjJMOpxxqy5ASHVuLfVdK/UU4S
NGKf63Rq08IZwKDu4n5wmP0eD/zpD3JgXuMHHJw4DyAdsxyFFXJ0RBOQHjgBSwEz
1YMR07BdPj9eXIsonkUTWNIqeG83epEyTDyCH4ZRB8draW48yxgWDArLUfW2BKz4
hi4y1V3dokA8p/bTQI0dR2ZozSsvxqDzB98sCWzzvXnGWMPj4zLGJOR5wwYk/S7j
maDO0Ys9PwjkFWNHAP7fLE8jrsYuoBXyBECfMrzKuluTU+cl/CM6/hl3hkI3tuPl
Vy95jhXv0Dtfp+cf6wLtW1Uv/5czykbo7qWUyGNrAB0IktFfsT/Or6V4MAAJ5Nur
NoIZfi6wPxcW1kwrKJNLHqFQwETerqJ8iG2ycJMlGFul8PoeixZBALa3VX2sL7PM
f/HWjjW+UciqlwW3OS6r8me9LdbPrwhnmes+ocx+pKeH2KBHjmcTx+jlCFBSz4wG
rARJCdREtwGEPlBmIscVyZBKegvhD3sm6SI9WcBsc2wTkBg1MUWUVCiKEIqpxX8B
aLuG1ptYJE8rliyABh41Fi1g9cR2qNE0UnCNqk54eHw4sYM6fMpFZQX6tbHJ8qjl
9cNknL2l5o5In/7V5XdOyPv7zpS8XYT7U0qidE5NCi4VxmSJMYHXhD1hgwfhn9qK
duIBL0iSZP6/cXtEBP7lR8b0LNYYtkeqW2cUMtw8fILplh3/VPxbSG+jCXSH/HTu
YFidOTgeuHMUx9hZYLyvVXK4oVTG3C2bcwDEPMrAQIYftcHvMu3hT7joAzV3B3YE
V8ZpcJB1eJQwRPQoHRBDoTUIE0+27lQbCQZKO67AC6wZl4SDAw03A++mOs+DiFE+
8K8u9IJA5+l5uOcFTHpr/D8U1o9kISM5KJ3JryvUr2PR0nIUIOxkWAUco++5KRls
UGDf+FcbnlGIw0gw9wTz1RDvGQIepQfVlDEgj8PxSdmgAnICbgPp9tTLTO8sXAIG
U6d/QpjUuXyB9rwQARZMXtzMwm5qqgw1feR6fWcUmfe7FV8OeKHsbOEVr2b9G08J
Xop93F1Yo8gjYUMJR9kk4oGWWXVcK0kixUBVLxZWsr8CVuun24iuvLMCGOhrPQHC
sulG4NTwALYwPUBODRMOu5V6Lug9RwbWa3ElqAO2H4Rb2G001kvRcQVdPJcJVlEH
qG5E1bRDoKvvcQhn9hEApzFRSAQ/GbEAIT+C8OhNSdrBMLKZVLrPRZKI75HSYeIK
nE8G6kdxgWjiugG80UCx6bir+9AWOdJsoWPTUBp6am7rz/fryb/xmhUjfNX1QWgm
dn+5Mi7YJ0AvEgc3/fK6O9G3XzbeSv/6bDlnQ6jq6OHp/q2LCrlfDzoItsgSeToP
Fzcnstziyi+ppeVH2HRoM6VpdzJ+eiRs7n1dJEDvYXEZFgehlgAHCcWo8NIGdyOH
SxT7Avg3ubDk+/D3MXSmjPdrYIVe+jwYkIdNq497dwT9akOtcqYXi5VmlkXKGoax
24Bj5ULtPKs2N50TeUE5fK+N4cpF0caAPLv0bIe29MxF97WzJxgLX2qc12WBGsb8
yKookZB/WdkQRvTqxnSbznVgpQ5wEE3It7yS3BzJZUAFe1JUCFg2uNmTUJbzuv68
LArd5uU0ORgDzbJzpNlw4Rjko2c2D3F5igoVwrQ+yYSAvydXsaBXQUjd+U1DyDKF
ICbNeuov8UX7GNVwTfTLrR3OfSHbJg9+UVJqvJMl+tLKLvgLifgfT1FH//+Pg/o8
Is91qcx29n3o3G9WMgEgjYQqWpIeGru35wWQtWBAwRoJDO0x/yaL7A/GGKT2IRMN
bQdM1na3hCL2pNjQcuJASNwmaBft2JI2k9GdtV9YGTP4y4Ultu2vgiWYyIeguoZF
WPTXL3e5YnT8MCCCq7x8Y62ockU1Yp/UtddkVb8mQeDs4RcdcPwLa7sZmMvEi+WR
nPVx2B53/qYSyD5NyysqShvBzanVgFHzmiHu7wUE5sggTpL/8FfFWf8ii4va0EKP
UWwll9IHg4kUaP5UAr1flnulJ80zsxtLUqXvxpPGD4VIWFnZUEN9Y2h9NCKSGOba
tBt5i2lKfEdbqtzPjYzPvb6zRDc1JmhiNQREDkpyHnvkCo7Yw9urLgLqXh/5wkcs
rt57OHmeraTdAD18MUxTZIFZ4AlsCudYtHJYhUWGIicNH5FHZ8wN1rY/K90kFaPy
II87/rwZrw4RhC+W3DQFFDDR0c+YQSCI5qfT1lBywVfeIBtbSbxaaxKRuyxIVPw8
DGJBioLFjEYZyvprL/1Mnc3XzfApy9kKc3iG0RdEN0pHyxal++ZVz4TP6LKiU2dS
I/ucREtAD8YoUEYBLARVN1Edk0KlCyFZUg5FMHeP6NRw9ceMNEGhxbNocJ5ccj1F
iLV9DPNfMxUV02n0Cirs3+xc9CEdY/gg6d9kolXcsGX4zhHDQ/EmvpVQyjxYF+7M
JtQ3XuBfCNjrvQLN3P+5wCe0qVRNrQ3HQw1vvH+SeTH7Qu+4D1EP5OT/syoBqGTj
Okq6i9HmKKTutaZY6fcnNZK9jwxBRdkIGh7CIcaUc6uXG2jIC7xx52BMwpT04rCs
QvemMBbRk5JR8YP8St6ygBz2a291HSQaoC60W5RNSlE723qjIuoQn1AdlYNHiy2y
pIPAobnt7vM9bLv+ae6hUMsRE0Mk2kOey/Fp6b+IpBPVsJZUOiLYkHoTQjx8jgJe
Sp3XjHpe1WPeDv6HCFV2L8CWfgM5nSburKcGshtDGkpPHiyvZDBtTt8ZEye/6bH1
ZzUG9ZvIBIW/QwqSs/imgBxipJaQ9Qoc+yUQZ/e8jaAeAHsfBJmzmO9zvUk31xAB
0IuEQgs2YSxXjRQyLtXtQ226nNtwQXe1dI0Flmj1nsmE2WgsRtNhvvCjCZfZChA/
7J08bDVZrxsf5E9Ztm3vY/BGCDFiayTSbCQ791y119lBVjTL9E4N5PQ4lJV92Vce
/bjyCG3Mrolym7qgAKZXL5t5Cwgvt5bFHXW/V5nS8bp+6dkIzQoBqJckzvGxw1d0
hUJ129Ys7wFrG5RymodlQRefcCTcMxwzK1fLZLlKJKjWtMEgpxxJ/JLEBHZXK/fn
Qik/pKE+3xrJtBPbc6dmwf8k+oEeE2omIH58lRFExek3//Kw8YT/D2Do7k7sfRPA
jTChpmpGrf0umDAih27GmGk/DSlCY+5tgjvjM7vwCD6Ms2ZaLbu1wTJHfcZ0yxQs
ye8sFwSq7m1dcARMf7KAy9y5e0gou4lAH1hELPhX3TfGca1wCEXL7EOY8aXSKjW+
jj9tZYfVW8FhzH3vlMjWE7/v6tFu62XHA+0hJR7Qu1/wuZL6eRBe4bGEayq+7868
IKuD/n4bqve8PEF/1mw3St7NxqrU26hql7f7h+OehZgXQ610u6gJqHWBgZ03gvup
KiGuoqvUZ3EbQSsy95UFQmUyaZ5qnd5Sy8L2Q/pCxEdS2ETsFBbWKvJylpi8xpXY
niczw4DhZYe7CSA+NTm2fR2Q8R1vIw2IqCyACtGb0h6CD5+tpTO7CUyR6H8FRql5
19ZqInqkWVL4hYjMzZkADYm+a7Pu/fvl+MQ24uGrwsixi8/dcFs0MfqWUod3a2yT
x6FkdOOwVhfhMrrXNGB2St2KFW1HEEzDbyIhWAsn54rye1DsPSgnLvEEcnTZNVsu
B2zn8MQMYvaX1AExBKGWFL+0H6eegU/xlFcF1DkZRQfvQdo61GSJIyl/KtAeZIgA
NMyp4nb9/hc2kT51Ustq3S8nHFK6xbLrA3d9KMhzP24akQ1AFqFBdC8H+5jiillY
ZlsaQGCxp1QXQBf/EHwja9gHA3WNF8gvIxPoD5xjGerm3aeAofOxZ+9JMn/VrxWE
eFvPR892dcYxNkTXhOtjvfs3Iywk9Z5d2Wrja5GsePQAXj8K8Z7KelQmUGhTjuzi
a0iht7RJNV0I1rNV/eWiLRxlGvzUXAySnbilY9RJgcat4vgzSO2Mc6W6nJoQKwZH
jUaGONRHvDiMVL49ASPzYjI2d3b9I85Z4CfG5B3MiAQg2fENolwaGdwmMr9QCHrH
OlZRq+y/NyPIancG8z4Rrv2dMbxIdbwLRMuQquNeo/bU74WX8BzheMbcgJo++h29
IkNlBiOemBltVLCV5/7pepGyCMQnG2nq6YyQfOOVAypHpPzGv2LCKEMmt8FPKIff
7TB0bnfx6nmnSK0Y1o+4amf2NTBTFWw8Mb3Rp3kHX7imp3mWbVwFPstv+MBpJsLg
f1w107egT2kpBdkcgDQ9eTmrh4uI3dUz9PQtyz2T7Nrf/0fm/eFgYLHS97n8kuFK
aqi9dyOxJgaYAnQJGryQ5zku2jhOZmeXhVyPaV6LGPTfGmDjOR8oUjIK3+J/Vy97
v3KDME+IT9nUPVG2geCNuDeY+YTyvzUZaq8Hdz3TcCXUo76EatZDEVrWq4+rePIf
sD1rAMFhVloENFNejZtOGeKoE8/KxiH/3gm0v5uDxIbt0RBCcVwPpwdFctOsjnWh
yXlK6MPLnG9hbyXjmmCLGWOUrscUnsvBFmrMKw2weZMSvpR8TodRjBeFWNJNmAz7
13DIeFUWYY6B6lcBr7P4TlG3W49diEtsMbDhNx9tGTSGZ8peP3SgVd8qWEiJT7HQ
3dochFOYHs7JiTbouwu0ZF/1dxKoi7lIdKCUw8dXUf6yxw0CnNNSsazdc7RxH/cw
S9akNeGpf31EP3tUw+dWVV4NUPbwRbtUx853hT3KGFFYyFl5HMEGWm6mpcZ1GG82
QG1dwEGVP1RA84sbbZItAutpKHnbc5uZInDOsM9MA5xkHQr4LYsOzsnK8rvSOHAr
n3eHbW9KwuoP0wr5TC3lP+gA9xPdyCZZsG2NNCgBUIP/F8CAye19DVWTfUBGVPzV
T/HlemtqUOwnHKTAAwTmMiGnLQ6TuE11rCo4nub966YFew95aCo5y41zZQvqDB8H
LBBhrWrZPsXgSHY48+EsexXKLef71CxWOhedBz/ReajuaRIB4VVvF/hpGJsABC8e
eSt+FHxy68Z44evxjsGbzMAQCGICNRviemGPUxbjDEmbpMS1wBkbEBvuofUeG+Ob
bcy4EpL77seLy7phHStba1wCy6HYUxhAtRx+ZoNyiQ/eovIE+BzXOmSukrc03uIM
myWh4zfUjMit3J9VDhsZoDiOF7TXu+QVaesAB5Ls3wGDoO9p8x//nCL2HlCzP+Ph
kTqNMr/altqymmNB0iorTLyiqN6AKqXyeQ3vhrnCOM0K7wzImKGWVX2DlQSsJ7th
OURzttgmfgnjB1QgLLzf/fZK2c1enV9xZX86Pjf/nPfs/LA70vRSbdof1lNegJt0
sNRLbwq+PWIp4axnNSHgr+Gt/pac9sQ5zWExMu64Y8BnGwlDVkj18Hjqxo0g21kl
luSupfWwnZ4vE3T2ZkhOXHmIYd0sWd7hjkAKlbdlsZkO962t7vLu89WxHV3lK4Mt
IeEeP7TnTqoY/cp6yuUBjU9i85LF7I+KAx402JXIL56Q58aS6qL+g4AvBE1qtCuf
hR3j+tyvIWdPoYEZfKAxxDKkkPKp80zea8u1RMBMBwMY/nl8y9aNUCqhtAw2Wuwd
yNBxXXitBv/FXfnKTvjNpLs0nv0YleEKaCJjHqit5ew7rtXANo2w7OVAArnGk3/y
oPYBqGcw2LdzAAxMhzVPPzj1/DutUT+BMqBlBzpaYtmFLqIeM2uy89JzdYUu+zXz
gayeopqpbL3WSkNgKXNxrn20U0q6IcmPiDCdoIErhjatr3KWDEs4Y+8RloB6MnPs
swcRs/pNijDVxbVdosqhbVx6fnPIJb19Krjoi9R9NkJF/UOGRIi5mDplCg/jOuC5
VA1T7Uzcotou6ul0ngfVHa/i7zTKDT64oTQMqqx5SBO0y5sa0asf8lUjB121IQl2
s+HIS8/eDf+QKpyNMYHZbzK+KC8RpJ8oYuR1A/LrxAbxC0kdTSxa7mmzKAVzYYs9
vHFtn7SsbPBAk8a3m0dU9PHsJM0F88EfpaiHrgi2yA9I5iO69sC3MyK6voG0Zten
YJR9d/AK+I3OohESw7kIVqvoH8HIDGtA64v6+yon2G7/p1jFG9GV3qeaYUgtV7gG
eE8w5AxG1eDWP311KAJu4T4ZkFSsCo5kS5uXcMiecBNdodK9WfNXq9uB7StV7VXo
8Yz04ncFQDcimQoKOaIqcgIIBmB7Cg5GDjGLF/Ezeb6r8lbFLdb4TEx+xeIuNXAr
PIb1p5fLILP/4ggH1kPJD3JdHCxW0XP4Z8f+KNwUmhv2+I06inp2rJHlxORAKg90
LierzOIvsUfAI8l9ENivSRK6rhY6VC5LROiyM4v85oaQXbqNL1FO5ZaP3+cUG7sa
bA9J8XVL+PUPUcnE3pRiP7hvsaG57eUrzE7fYQriZOE1A3IPkQ6yBqS945JhSwVt
r0wTBnLYd5RXxcpA0iktjiKjLrWnde8/6WpXmpueezdkaYhYgQSJuj30iXpdOSm/
XGyPoNIlc1bKwXBFkmSjGkFFF4LXVB4ZQNe1ZZI0yW/6G7ykxYlbahv4+RlB5qfT
DWmw6kl0T2dk7Enk2U+aQ6pdKvSWut71CBPRtO1im8uesUUzBQXB4Ryte12tcvLf
J6DTHOElswqV+i8dRl/bipDtl/QuQI5ZkuxgKD/L/fXEuy2fCdyo5ObUQoE6qNjg
aY/ueqkjZsOEj+Ak/R8ZnPC5ZZkLM01EquRltCQXx/FE6+Q9mfkfmrPJmkVCvxZw
FVPkyg5ECAmq7cNYC4m9FNwoM/V51ANkFJJX/UsDNuYZ4azNG+ffQNTP8BfS4b+u
GQjeULlurB7lFAwjE0vxUgx4V3xUssTvVoJa8dKVM+PlZ36VCPzkTdbyiF9hsstT
+e1nw2RTbZquHNbGxz4i1hXbl3IUtzkYOlqa21QJCzkcOpS5l4AFlvcL4fQLg1q4
ax7pt3E2BSgtlUmJx7h6acFwpEN0COhaMd5Q0lkHftNk16NAgkIGcH6x3aKrH36T
e6WQjoAuZ/+1HE8MZLC3daNs1bNoMA8xIlxRKdFwTbmD8+7wp1BZx9cYUzWAZrM8
e2IC1udyp7vNaLAGsxh4+s5TV5W4cM2USRPkk98TJm7AjRICOF5GmbdbJYVKWH5G
2c60hBAV7U97ORa4GjCZXWHrdPUzSGW2eyzFz6bqdR8CUDiwEuAWWroXMkTQc3aH
fD51AdYmhEAaZSNNvOUG6GGLMXlTWxHnzD3lT/E05IexYmcCpcZVbI16IVvKKKEJ
gMt2l2jFhKDhlvEtf3LaL5ADSOWBXhNsCuZ7iA3tZ6c04Krl//JOgchHdY7bwd/Z
GyHF1zl0tkM3Zr2Bx0rALz6qM0i4+rqEleYnpZXZeitCzbyurEfaRgNMW/qgArU1
bvwdCxZaoqbVxS69+zmh5883eIMtjTl/nSXZPfBT8/cs/bE8bJirNag2btPpZb9r
O3PYbTqPJ7AS7CE6pC9EoAE/rvByU3WQRGy7R9PN3ryD6x/N8DqLcvArJNIvCifR
GgSbkS9x3etFHgMm9qDU8A5ivvsFt6uYQrZAWirkYqOsIZ9e1A62X82CQlNcQl4n
qaEQyEcXEROaxbHC6uPGCjsPivjJ+OYHpVCG2t53uhVh+OSC8v/ci1Pj9h+rLHS7
HvCN0y2yYLLN1KB1YCItZrsuW4vvCUxGbXAdUabFZxUztQwFs9wf7yu8bJDol64j
slGo7eCKqNNH3OGYFDCSsYqyblN2h9AB94ae99e0LQjnGiby08WaV39HRX0cRJWO
1NHhZUVMe4qOReSk56MA679Ec6EGBK7sRnx7lBBqP9Jj6FU5ilQkwpqAplDzSV44
q4TliUmqlFu48mJeYmnEpEyLY/MOBaOSb7cIG9qUPj5ItXKfZWnRqtwI4+AbM12i
Vg3NiHibP5sHcM8t4GZpy494Fy7w8Y4Gemq5Z5G6WnRchUbkPmnudn/tCt9Ng9lx
goQ7ddIOdBgTieN+iZ5VdN5u62XF8WLhwAfRqcC7OlbNB4Og29HflVirHWM6hMfh
1o7qxOxSOeDaY3ByMJQCoHdHwzmVhNqUJwk/LArg6XsshzF84FZY2Imw8NWF+hlc
VVRx2bAKJPCp4TDzdHrYaszwigOju+JiR4ArURJrkZYAmt/fVHiNZDlHqc0Wg9fg
K7fa829RLfBe95LMpEkpr297jGsq/J/1ExQICQ75lCjUipxB+Oq9eT4lJYzHa2hx
vlkLAbbuVvdA0iOFbF0FpVPKZ6FN9aswHf8zjLNomxOw642kHOLe9Aa09TT/64aT
ZmpS9D1aSIbljLVyny1ckNDyO0VOSCfsZeLrd2bfETdov/KOM1UdGHquum0d/ih4
ERWBZ/3zBGburQ6m2vHsdj8zQbYgtvXo6YBo6U/1pDNvKcesxCHbyT1Ha1bsPL6L
Dl6L0t69i13vHtKhCsB9+SfTKNWdI/K/4LLCy/oefMaLYqeOgRPKaFgBgzfnWY2B
haYnP4bcoxsGTsq4S1n1Alt76TOhQcWGSM1797YnjfFTDAgPWHjOR/Ooh+YqEmVL
4tG2hjFaBCjEmuaRb5+PNOmsJT7xvis9WxP820QYtacqBM8y95dQcV9noXq3NMJm
jzkUSyozK6E+gJb4Kqcga4ujwSa2+1AvKL1++xPqQ0ZhiaBYVzN6m9M5PhaCESOV
BuZHVqtZIJSgaoA5/NOufuoo4IY0fD1yZkeyiOEIGHDb5BCBVhoid3IO2suW5JfD
jDLQOWIBhSHv+TLh5EnzbX0Y2o3NpSZiddhqQrofAygG33SxXNGhB/m/v9L2BYUw
aQTHD0e7v+MXgh+6IyLwrEot0CieghWfUZQDxZwBRG91u3zlMVRLfpRqdbTCqUpR
a+QX82Xu0J2kVQrKKlZFPzdHzveyO2rt7I5jnIspfjUrM7k/qbx9p4AH9COyQlJV
aOt1RqoI2bQRZ3/a1Vu52iRgCNy6qMprAr0xkDVezFsm7u1uIjxYqwLsM+qaGueo
mWkXRWKTQscSUuWs/zyR4wOwqb9CULm8hSN8Neg55i/tnCw3DE87tPrwyraoY6Yl
6nBWjExMcPZn4lI/Ipf9xbYNGmI8O5ypBgbpXlipbEeBO4c5uirL9Z051fPdj4l3
Wv5OVepisRfzlNZgy/3b1m8L9GWecuLuiJNuR/wN9zQWSfKUUi8Nsz9jzv0k9HdZ
iWtj7UckRxc3N3FdfR31HhzXcdPUyAs2bxdPBBXr77L3yGQ89/F3z95WYVbCc+y/
3wIQLTiO0rpEathwNTlVyqDZSoP4568LZKr7k/JmO6hJfd31JrjbPFfORX5CCVPE
4i+MsgUhMOiRR4HzUJmivR860IV52TgAFG5k9MZnZPPdshLXDGuBMR1eOIwDE7GU
2XDhjkVBdU4cj0n4hQCZVsqhOT9apj3OfFrpLlYdEnVYP67B96KhUpIOE7YLD2Ct
88rfuvypIvmdoxv85/V8eP5u8oLOdX9g7W38z+qpgavzvQeMqityah+Hwbp4PUWH
vWRwT8SgW+VH2gPisbXv0ghTdiGj3GbvoaJVELqiRAUaxvcesrh7fZUrLh43siO6
aQbJXXSdWQs7JZz4YX+6gSHZCb9AwT09WZwQUWPkdaOgT0v5Xc+DIazcbkrnSsGz
Hoe5qRaA2ATNivjx8P4TxbzF8QD0zWZw2JSa/mrX2eojkbQbO4Y0ID2xkNC7xEhl
f1o+A7m3vOhQcsmYRXqgTfBbii1eflr7ryUKCHQspJv3IHUInzRDMBiugs9sw0Nn
RdW6rMWdvKZSbJy3aHfwoRSd802LoS4+9LXsigtG4CJAiIt8n+Vqpn4dcbkDAHO7
wiEm1X/4eOn+PvBB0WEG7yIlrlTtfBwJrUZi9dXbRNc8AhaC74f/+6u8k7y6KOt1
aPSu9HyYxNp+mdlWhtTQPWgfsYwk2zYqdw1y6M2KDVOrmPoTknWXns1tW3vzhGiD
4efLdLLFgT1+5J+eC6onEoCcERJ11A5SrVx1HDGrjTyHNb2PaRdFnrxpbT9I79Cf
frTZCvoFFuteFZYvH/ENTO8r6dNDDnmvvE/mzxEjirrSE1PDZKTTlUJaZW7q36GF
+KQ5p+uET3qzDU7Aiho3NOLeXMEDekcMMJXddfC9Q92EdZovQpkYilKoVb4PjHHC
S6XVT9W/J1lAiRalsATdTck5lEX/kq3Wj2Lz2kx1CSJVkyyCHBhgkuoBeDSK0vga
EQu7gz6fCHbkzwoNYfPLhGfPOczePHcpQVfu/xQVU2rM+ONxecC2Y6JSdXWJDTR7
i7H8Ok2pH30EJNf6w96yj9G6TnC3nhks7ph1vyXqHXG4GKPd8zqg/hUdzzaVvnbX
NyHhWKHd2NiWBHnjMxEXyoX4QFnThvwrCRj58LJ/l7Crz9dzC+wVc8FVCNyBhggA
x2fQ158Q3J3dOCywS2p9McFHgfBiKkIyfiuam1wnkCW5xnZeyxWj3VnkuOvyMHFB
lL13oAC9m19wGfdWNE67ywuTw4TySx3nTYqXaliGTKehBgYo7tQICT7xhM7VYtRL
qhdZ9HPv7rz6eZARtXxSnRq+GztYtNWuFtUITwOIvFDeTPBGMllxAYLaGBe5HWMA
yqkQCJ87l2tEEpJcJ8t3sirU/Bt6H3i2K7KZLbeO/1GLAfm7c2dRSFLHukFsIW01
QiIGrI3rHsm7IAYrqS33sw+bTybCdvSmIa/sGbUwtuUwKwwPQTxFjTcSdPVWr0Xh
bSl5h9y6AdWRQM5t/nsmF1l0HjhUxlomw0xB58I34glS4l2plGsewWveCM5xX0sx
dJTr2XTPdo8Zj0/oFGWRemKOzmk5UaNeX6Y5dc2SSCbRTkp7cS4623DxtWXPm8Mg
xSJihgj2HktdAo9060Zx0nCkOO5qDcli13kGhsVuIRBG17z4fQ8hgCMWEgZ1yYJ0
NU6AM2Cvtpr13bAwaC+6Si8QukhlIUnmo2/ne5gYXiSBSFCkBDYsHT1Df4I+w59U
giF3ZJ5sTjmTa/diHKc26T7leca4wGuxNakpVGUyh75o41/f82+RygQ0FuFe/2WT
wBaX69RBLyHfods4H77gN+0Mo8Cd2+BQxABQhR5hkVpD1R+U5SFao15bUG/DGg7I
eBvnDBV5ketcbgvKe8LGBViinN00eBNgKmPh2jwee/bybSZNJB1/pz4yRX9WV8R8
mkyL7hJmpVtcE3Hwf4JZ7L7yAEH++aAP2cit0QMNfXmExilJvxOgG2ANdGX5hxp6
kg3DYWHnaHupYUGxGIN4epwvRs9FWHBZHlzaFfvHo0+d/TKwwpGB3YWhve1i7YPa
Yg2gUlVP4nFaNKIYLPvJoM5PfYloMKHblcxlykYJ62QgTXFaTH5eoeFG3F2l1haE
3L5uL5lTTxRxdIHfYlydIcZpCEgQp0f4OwQ2PdWnuwyOTlTKMc7ndGgYWdbHOt+1
0b5VNnsp55UFp0DbXUdDY5a4gpUBNs68jRKXQ0jZW1e5vw4A0Sz+erSA+S/7OcIH
ddmJ05bhfOytE/kq4EOGExjL3FjIFT/xNhtajCtEMiX6qQo0vQ2nNsx9icRjc/oG
qaAa+ZKZknqK2H1AtIxOTgHMBQh0GotHkFswgTf/5g52JcDIucT0GgakNAkNY62E
GtTFY1fbAERrujjY/2ioMtm+yn55S1NT7CCpOYvPIxGxJ5u1xlQztEWTLCqXfVyX
BqHWMAKQ92X8K7EjCfwQP6in7bORHGfwbVFa5i2NvzwYo0WcAOTa5clLC1Ed2yuj
yew8WTiCcgQJWGGZo7Bp0NrLaJ1lar0KvNvp53ADB0G7ct3Xo8jTb020jYiCW/GQ
CNV3a5zHS+PmHh0ZKywwqQVjnWswLmYn99lx6RFHvvZBOgloTzkA7ZWVxuLLA7Qi
eVeNGwnyYqeZM72IjcKyT3l6vJMdpkX3ntmOlTTfJsyg/oTI1VzFehwZUI7YUOfT
1HXVcsMrmzoqCitDgXsPPLIQhUSqxN4n056XCud4NoXqGG1s06xVp6Dtu732l5gF
2E/aW+Zxk93eRk6d/+Gdp0acguXjbowiSV2ujhoR4xa30cZgFUQZltOKE1nHAY8d
A6e1AfiCj0F+8EQzqBBVrLAec5kwsIi2I+r/+jiEniFJgJ+k3hnCdLweaIBSKG//
S2v9M8Utt7LZdHL08QNT3iw5KnTVGvf6ybfXSpJKQ5U2EVf6Vb7jRzFsxd12rGhQ
wH+VsOKZJcePtaf3oHnchOtNXXtIl5aJs5ugxysKqJnBkm/L9xLn35jqybLG8fRL
tnv/M/0c4hUDNHyCrlaQDsciTgvL46Q0eM5sxOXgTKW0EyrzAi3yz+Cs12Y20vtI
QuHOwZ6WO7LarqGLb3Is9Svc1TXA7yoyjJgi+cHRt4c16a3X3OzAqCssE2peWt6B
LZOLGGyFbhO7ePSlpk2Av4fBoCmbnav3B7BOdfPNQknb7Xha3RzgN92e1orC5piu
3OyXzKa3PPTJD/M+m09NZBRcvojfQPCodiTg0RWKzppC7hqlz8Em8koZXRJmKxzk
Mpvm4zLsY2VqBepJMCYTUoWIeSAlmZqBaXkj9MVBb+7dKDHNGgWxLduEycA9Kem8
spstT6yIdMuptA+JITfbWMuX5wIKvkGZyG0T2sZaxs8jSfJZJPLNrxnPVZaOY56M
lnIiedma6MdZCE/wrSy8Pi9D/rfoCy2AUjujPg1L0HgBuoccDvtOiND24/aWkm9+
QrBewZISPmEvD6IT9wPT8ij3oto4c2Z2d2Y/kBZJiXmPE2PSm2yUOsezPzC0Gnfm
ydFQYmnDWqtOd6iKYHerrbyeHHgh0zpATOdQz7UdK/U8F8JPwHmelJi1+4BH+h3q
OXnrlx17nm3fMlj803qU+xbPBFlEd1igFmgQjRIBMzfC2Qlu9lKArUe7ZrCUoR4P
/kdi+r7vg1EmIvJgERdzhnBRyadBOeBz3W0nPN6XhrcafigkBMLPerTzSxwRtW62
o6zYyucJB8y0GoxxOmxuTqLcqsLl2mgShQy0XLB0KYJ0MLvIenScvBkJ+IvMjV3E
u0TGFQ52X1kcMHeqlOH43t9iPJc1adtbP25U5shWnpBHVCsV5eBmK38WRTkyD/me
RN19eaid+KEo3TrugPyONpR8hD6CGe7gnN8SfwIKdMB81eBKmCG++vFLSpC0mTpS
3v5YsQjaBh2P2UmQ7XEtKU0/8pP+UCVJpAkC8PBCsbHWnVoyH4lu+6xvanv1YqDF
+wyrHyLpqJvhei9FX3mDtMaxWjk/U+eeebMG4rMg8JS0uuWdWMkTqAl1Jji27lzh
HlOHj6yjTV/WpqKNRpOH58RoJm4Cb1Jq3z8mujqjm5IrCrYdrfLD+MSolQS0c18n
jlkN6Dwz9bxLJ9LWlLiupFvFCq/XqxlAaleKDTP8nWPOl9LUWyppK6MWJg1j1BGK
qnz3PMq3GoKuT/W+r/95lek2z36DIX5dw8Os9/oqGTO6AQWHl7S2V71c9YfYQuOi
/3hcxfeRXTlfxRHlN+eDnZfuQden46tqYDtuC+QXg0vaxBvWExkHJHnyxJdkP9Oz
K1fnENrWuj2BeaPjeRDg7vuyx15Kz/lHtfqzqQj7DoH+O/+1Qbm3Q9RxaibeJ8M1
pRgKyGeNhEKdp1CjPjYBAIujZV5h6zYeqHBeID5ZIvGLZHahqV+VvleUuStVu+gL
KmJ5PTb/5cj8SK9IwXTajOkgSvxH4uV4wYgTSw/G2WspCbhG8k4M1jyDFnpPaCUX
KZLxW00oWLdMrJWKjMZuIttzW9WitLGHRLz7DIvqnqXIH+u3YOFuKBMMgyHHLl7A
dwMfkVAI+Omw/jNgNMYaQTkYtvxvZ4pglLPzOZh9WXs6pOJPNk1TRg3SDz/Mty24
5uSogVQXsbakpYN5jYpZI4Ol85NhHpOeQgZtJz2ybRAU+jH2jPjDpACsJMEHPDf8
32gKrcC9Ys5xS8mnULpaL6jZUk0TDqBQbqTs2icXSXHU9A33oV0+p96vzc0vMxN8
9RAgTH19fN5dOhpNQ6lED3ck/0UJeJX+G0c7tqE7QVJ615jYxVYp2YFGHrhUNJCw
WCn5jZy2xcrCqly97OnltaoUSC8E3Nj4/+rgHh36KgWS2KEh0f/3+47GjrbOijxe
Cag/Qm7D10Rl6eVXMKY6duq+LcEvrwdUKDXufiNuutClLATZBoQrrzgCWDW5NOEZ
bISlQpZ+EsT8Db3Tmoc8mggq00FfuSeAN8Ue5qF9jWltECni9W1Toh2Tq0/DQcRx
MR7Qw2taQt6Ou/awo/ZWW3tmrS1xOi0NV2+qjNZVGu3duDGflP8k8aMEozTqknZH
xW2JXVCxemest6CYVUPzYlD+xzAXgY8p6rffKbEOzJMw982irI4UXb6ahwuwiBJs
3JSz6jqUuCDhs0GT3wDoxXwF/pVoEji04zsoOMK31ceCsZVbdpD7S4tAX0FK2BgV
exOGLeFoK0ZCckeUgJbWFGWk1/ZvwMwjRl6B4CVjPIaxxRUgwiK1zHL6dVjD8G8p
nZpNgAlPAba5ZIQQkepS5QDkQ3OE1UIiDwp9jga+Ofz8CYM+s2tdxCn/6+lHRZdz
OPg+BkSNNhFT5QM4dw3r8BYYb4Pf+WVeQewJo5+O3rkjv41IEI2qkD3MnGl3RIO/
BfPBM1hqNyz+RlpFuFLHrG1DEfZK4WsAZjmuz0r6WqWmDvlF4cMRxn+2qd1pt6rF
ql8MdWFseFUU9hknemgpoZCSCOEG1bgAyxkLm/tCjS3TAn/S0+EwMtSNaE8mx5YM
8ICocO47Uo8OY4G/n72Bbcrl2z07Vq7RKlnVqY/89eIUEewY1PfK5wChO30xI0Vv
blekpwedGKCVi1aGihfWvloEmOKJQvhi3hrC5tK2MSKl8+NFxNO+8KU+fIWiiZXO
mf5zYpElFn1HKeJWKdsbV2Zaa6TNnz3LiQP7zAM83vhX2AKgp5Z/Hsg4pO1TgNQO
M0Q7BZ4z8WdFrAoTb+0ZKcz0cooIKe7YqwWnEB8TLmNr8biIg0z2DXQ9thp0mcae
iLudyJzjLwtaDjL0XpC0KElBvPo0Ytq9wU7xAqc1KbVJISK4W5hbUsuraFd2xi2R
2Rj3PFxsmCI3h2TpSHZHRfFDLbSODCXgLxrJVN+OGxlJoq7olpkIw/7YD8sIE6yE
M1+G4uBoJd4GDGCO1xsvi54ys2uPPcBFvBiVL3TlBErz6sXNKOAUUjV1ZtuOMs4G
B5tMZ5bKzlquWOco6xsohqUehn0PtxI6/Q9dDuCaEZXphCgYq8uXGGDDg8QGfyk3
N/TODO6D5XsuN3dT3Y5uNOfyEZHrXECbksAe7yLi5eFpXdPRhtoHis3zyksolAoj
Hv1AyEuC90qtdGN6jJQPEa9dJEd+mik23HIaATHd8jvVtvqMZ2dKifQ0y7SCa23v
VKCUeGquAWiq7rFNlQYzIwez/eDB1wQHRdzWeLTV8dLIXZ6vgoaNzmO40IpWiZKN
k0QoL+GlD8uW6o/ml81x2NFhbEAvcLB6HnM/eMdJ9FJi1CZZtQgpGx+1Gk98RuS3
pL2jvsNX+EK2h4rj+/Bu3XNaNq0MKkgxZ7UyzJw7SaL6mw/p4fXm3x7PvSPgZVBH
6jMOQSR1+0liUHOqJsgS6oXjPUZyvWMwvYryt3JINubjpVIFgyp24EMC8Xslg0uQ
M3IptoG3hBp5HlAN+D+xXkfRvb6lc1VIUC7u8ocLXklZ8Deqa0IsaXe66RQXSjv+
bmTwmDgKc62X9HbyXFyV7d3lvExyCkMC7JI2OuZbWHCsqfaVbAvMT9MDP40wlvRX
4KxWm5VxDrdFAzh0n4bQEVu5kxrBZilTKebJt0AU+whtuUhvhXNXGHTRQKiXXb5Z
4kvDxpM9rctPb5QdK5dDRXXNWdCreRmBLRipLW4FBCFDW3gVCr0t/vEGG5DQROgY
MYmhWO5N4qC2W6J8XxtKX1YXnYo9/bJF1yZ8LKfZEQ/dY/jyZFP7Nt1WpEi7jcsg
WZItTkLoLqyuqyB1XO6bWK2wfQYd9vZQAwABXt9MJ7Mw9NvtR2mgt1KhTLmc+xPy
EqgreCvFjutpGFbJg3Ix1fiah84PKxa13EbjhXoLWw3wFwsiPZtUvvwW0mbRxGBV
V/bGcuN8G+Y2xsTnz637eUZgX85jPYCiGmJyuvZSkR74tkx4ZyKgpmQ758WJMofm
MG3vlEjqRFexnHN0Q/AEbkCrkQRpuhD5UmaYa1sNt4z4KGPBX5UTZkmA4KxqFOPD
kESBSXYsMlR7yOsQ40vcsOyY/dTYpOF0nms18ne6oNjcJtzbKZn1VD5EGMRITwbk
OYqmbKAEtL8IEF4opReGpRECxXJszOzn/K7ORUmPWW0fq8w2Xi6Ylmuuf03JiF5n
mt0qrAGbFTaRXOHfzMoNzjwoiwVbQfMLDJ2wzQmeFMMdgkWp4szRfYD+91uKqXMp
F0LIa+bs0zjNVPi0YCJwAkXc5qTpwANy6g1kkOKvq1QunudZxsu+CEknZ7a9vtG1
uivn+Quk+MYrwo65YJ3ktTa6hLQNvRD1+QbtxGs2H8/1dF24aLnpwe3gKasK35CU
Inyv9UeuRN/KHazCmQ7i6yZAXF+/ZQlOtkgRCs8hZxtK3IMC83ZDotOxWPKWTIAL
OoLczmzZv6bnIrGFnsHgNQC/mf3Dnh5ySUGx7/xuNt2c7NlIRpDhjCgF3YKDx8mF
SOJTTVuP3V0IPArBNw96W2wwqR5VXI/cJc6xXsj703MNb4owiQAcnsgOddXVDkSg
zsNRmoGUnB1SZpuLmHZjhateWRBOhIkSgQKYEVKgVOtEAQC5p1bP1M2q/Mq6HTQb
58W1TnzeuvU3IgeN9c87wt8q4ZrCHrc0m1y6bGfcl8SuhOW9n+xa7uED/tBMKVeW
Aj7X0XrDjeosRjIjRXJBM/eX2Bcgz2lz0vR+wEcep5/4OXl0fEy1DyJFpK3xocz4
UfOQ2uXCSGaCsONljpEnM7J7jvJUmeZZfz8i4BVyzPQF6GUepTjjwce7Ie7NtXhO
Y+12ITPU6ii5nl3Vbx13PvhIqaTUA44YOepnKgtMXubbANOPY/C6zJgnwiFVDB55
9Pf5yh5pKzwHmSCVPbVIPK6Cq9ATGNRiHU4OoREn8q7vON0u6+3XJZDKZ+/PLdeN
uCLV/u1zQ7EFI0FDH2vw3jKOiCaJczOFpB1I1IvXYnBBPydLXIGz/aGRaMBcXGDa
NOSioL+Sn2OgyEzejRsX18wK3ZUC2tt4T+IwG1TH3WY1WlRQ0xOhsXgpXwoyOEg+
XBRFfYb2tR1Fle2bF5BBjV9pNhTVZfYs5bZYRi+M0gZqFx75ymxaGxJMkbVESRdY
mhCgbdjkAZnCP2wq71i4UUcVHKAvK81ZTPjy03f7TNS46ifqzCPQnB+yB2ribN4N
+LxkyKHxfu+CnOTPXTbv8viT86oKrQZ7rBQznF5JX5OF1UJEyU3aVT4+iP8HpBmK
ApcDBNxX/7Mr0CIFGU9UEScvc+q1A8E90aIVlkRTRRzQMXyXq391Y0Md67Mrd2hh
sYgJlloxFgaAlA/fNV6Ygk7liSLmFhMI/WqMAr3W69Fu1SOiAsWRWdyjVFi45D43
VZJqkTT1R3+rjkG2krMol3untVoBpdJw5P8LGe9vakp4WKERUtrKN3dg2p+Dkeip
IwHcVe+JZYZAAwTXUOXLP9LStVt4a60dHL6BsCAE4P205nq5vvRacjbbETuzmWrU
m8A3INw6clsyve5NhmhCAgVaEEZ2IQV2K9EVayt1jGGQjwkPxiSsBlDwprVYkPxA
1kFEF+wdCISWczLYzo/ugsMMo92FMbTh2sl/B1aVfRvz12rYnYCUUBB8vNpTILot
OZ0EbBE1fZ/kBt0DAL1Y+tbJxDD+FxqEMixAF9OnY0imOaub8o38h+Cr9zg2m+bt
/vcoXFxEYAJnQBx8LyP2yyx4lNLXuszsP5gItgdhiDqd5h6L2UYHb8SbYVBjeMMm
cE7MV9c984+lKiFpxn2548S0CWfNUOVeUJSAII2m9bGgedKv/N0x4K3wLYF/EUzk
FPvqGxV4YZ9cXMe/Xmn8szjL6TGRpVam/Ba03uLuyKbb+aF/9u0Bc53uRGnvSUnX
43ZtPCXiNhv7E9wnDNpR8QJV2S9MTaqT8hrs+Ay+RzKrj3yR5tXRVSPEeIO7OtMS
3niYn21NHu4b7a1F2l8pSrpCppJadJ7hOc0B3a5q5dCDkeK6nnYaaZhUM0k3v2B4
NDgVxWT20ZpQ2h41QbES0MyLcjP+cB8IlqQuHOLDhdRZjI2JfDzL4IL7fKgyzv//
XmnCqg2VCA068nw0eKfGXSqOy/o/czwURdusfeqYTgF5bUdMsQDXnYllc7XfoZqD
erPjYYAq9GNiraww6ybrxXYTiDbN+QdHNsOqLxkgJBq8DiOiamZxqFV/TDW87m/y
RxQqcci1zbOyKD7s/BDRpPmDgN+GqwRa6WGr+d20HSD0lQErWXsH6wwwLE45VSfP
YBcPY4rdUyUkN4sxWHKs3Z507P+dcB3YhdePu4R8e6ccrKTUH5A7LUGsCfqUCFZs
Lx3jNMkD4/OfgqqugGBU2BByZWrJwy3bqKty3K1/6tFH5znVp6HWSVQSiFmZ+tcf
PtlEQAMBz5zAIpHA568rbG90ftFx7/3UchE9I3kGJrGET5Cv/hMfsJqj54TpA/qQ
Ka4BK80MPDascsTnnLnWDhPNCV/aXgtqx61Wcgq6+AOycAGxV1AlKVCXwpTsDC1n
r7lvcVfhc0dLfpvVES+uL4SrZ+jyCoo7DHdUq+MnqsmrEwkiuOiTJ+dY3AK4tCP/
DBpGUvcxjdLipa8CnGyX4IGlyvu/L5V69aKWJGjmMaXYSs8vU1B5oecNC5SMXPkT
rse8t4Fe71oE8yEu2Rn7ccXD7lt3bdL2j/jhY8WfD5OTKNT/hvZ/E8BbdpGYX1Jj
Aj9S+txDP88gnauQ/FAzUJ3wBcpLI38oeaaCzVdUUQ3HZEqd/FFrwcCj0/euwcX6
qegGtaF9dIEzCJN2B/X03I/nfYVz803oY83zEqBmKShnZJ/fOuLBpiapM/TrcKPF
kH/RfWUka3JjDNDCnXzfrUOJ6/KBdOlkzw+QnDyvD9c2Sxz2twRGhrkCAKtP+dzf
b/gaQgTd9icMxCyIUj7iQdvleuA9hhj5Ij+HS1kN9XxCx7dWqAyOect6MnWx2Dve
E21Zqr/g2KcEkJnldqaS9wqHWEoBCIh4VbTjPzG8necTWO6lmGeBwHReeZBfju4K
ia0YTVepyrspERXXyKuKKJrkA9Cd5jCwkY2+z1rrVYiNEdn+c5H6yxao9N7jIpSe
pV3tB/vx+5i2y5VIYKyoUNaKBNsStZvRhOvyCzq8iBZJOhGC1TcoaXycP9bGjs38
kvdLm2hFl57xZvbCLuL2zMQqIRhUfGL1zmyeZpWkN4AndOT7d/nsq8JDhHqT0yqw
G3xkj+EcB0dbnX29FwiYIMfbPeI/00X+NK9VJSmsJCMCA+l3mCXKeWWm4vZzCMcW
ytEdVhht94jSUKi0tya5m+AfgZbh4SOPG4iiQ+QVUjdxjRuRTbLyINMG4lHVU55q
cj4wBjMHhqE4viYTY2FBfHRvJSpMgNC5oj/u9dTFJc4vyYAqBDLJldn3Z5GMckEC
y9yxHmnBrJMA19DSd6EVAObAxobFHMoqa2aiPRtZWiCgb62z/2znx1mIP+EyF7S/
wZVKtX3V8/gDC1X7EUTqV/Zgb4csGqcu15NlJ6OMvFZfZANhez4l3QaSa9IXY685
37m9UEsmOef+nAEPt827yKP8IcMqa4b7JbdV+di12ltQ92YPV6MYrkylN9bKZIto
noy69CKxkUIQRkrSHdQ6i8bga37CEt/Hg82IYl4vGrYTGwNgR/L/acyMvE0wmOu/
x0Dov11/36Ua1lWNJbA9a85xw70iVEhCsjWqmM4Kx6t+wF1L4HVSwH/Fb8O4evL4
SwlYN3tdVqPJ9EjcMZQEIKmFM5yR8E76C50F7EdgV5fIIJ61d9+FLFYQuefA8nhS
zW9q7aZwJitwAJXaUd41k5W+NFmhLuzXFYrMc/oDcRpPy5FYZLMsTHtuxjI1NnOx
FykxqoGStZrPp0LaSvfa/J9aw2ZCoiMiRiRP4ycnnM/9a+30zzBvllkpeRu0Gl7f
nyizjxnaF9cR75/tcVGes8duP5qOeQID4WgG5EHJMy/YnPACnRyqqp9E3XBEgjL+
Bgl9tL9fXmCpzQQCuYfvA2VNK5Fd8exprmAMxvpefkzxJ4myCyywifLWj6I1rZ2V
2w9PbKPBy2jWgKTUrhebqeB0Z+LXd2qxudOBhaOc83Fw+/kDd+vG5zVAFFxJSlwT
oWPZaS9hxp+RFVLopt+3gZYbCQ8GezuNxkY9IhUZ9uai5cuDhIS+Y6E1qgwcNkcc
Bs5YffaCzVjPY5p8duyWBt7sGQFcOfOZHDm7RBWS3wnXzFQx7BaONPeehUGgEMGr
HWkeKYAAuFNt0LtgHDzs7xRuq4bTBZvhOg3ewl01W0xtSk9L0tcRU6h2UgPolwsN
ed0sgOwNP0vYxQJeCNbzLzDXa3oCHQK90MQyfHBPBc5dfL/UU/ndt8C+xsqEAgAN
MUseOljN6032vHsPZNF5XBism6orNlDOlz9NM+XZCXfTWh6S4fAKcnK/ylm/EFKS
MkZjgoo+aEm0rnMDZgsTcRTe1fLwAnwTVZdSiFO+3JP9pErg6wJIiXEEYXnKGc79
dPdsbctSgR6KHieBJMEQn4d0zZGWjezV3taIM1zulF8IZUtsnLAzHfOVZoT99Szc
QzQH+xuSvZEJKyddTojwuVq3D5eQLcJG5ggd1ihqB8W0j6iQMuciaQlIVKWRlfnN
Mu4dzz8B1PwVNm8SDPAvEqg9lSmD5OJBvcvm9+tAYlUlo5w0tAUfSIsV4rH2G6KS
IbgsnJRatGQED8ZkRA05fLFqYTr9pBPQu+lLd6brji3grDEZJsGj3ss4lCUhDRNj
aa4/NXC5zXzJXhjU+XzKFW29WXAoohg5PKtpyeEPmSgnb5RWy/QcPEBfgaULV/2I
bE2mw90xRSpDw3QV2ybspbq4tMRFGsE2rM83z/U8S5yCb5RpJCVpSB0T/icJ5Ndj
ny50VG1Bp+mxcEtmMdVVksc00PxPnW841rV0gWUWSCIyydr0MaoXiCIIDGiAT35P
r1kloqAbsVIP+rofu2qJKObecwO0ilaV9Rx1bLEKRCgsOoMswavM4u8m0A/05uFM
/Owso60IdV2KLAFaHNZMOtXQkawFEGnmzMKNGuD0WcqKhebvDOaM9AlMUVjFMQgS
YpmUGv9RDVfQyZ5mlUjCaN31X9Ap5cH6XgYBZtvzqzAHFbgMhjSWVNK41VxH+OnZ
pvMfJJf7iDI+FcKSYTnQO3oUdG+TAnl4uhdm8PHu5IeD2St+60UYpq8+D73+zEeD
FAfIDZPVM2EPEmnLzoKwxtVpriUlRgICe82XLNfLiA1C4k7ixMGbing6fwlGak7f
W0Dco3URVgmdyQR9x7mHqYncsrYQxJ5bcXeP5Yw0mJJQZjVkGBjxkvfEcWY2E5pI
l34S3NT+6cmg8EjM/o4qdylm++7kILUUFLtpAMIN4KAGQY6BW/HxQEmI/ayWfeGK
c3uDtNPouRnclpMbOoTeh5IzemCaJM7gS6oGMGSvpdqc8uUbTLCXs3joPHRy4IMQ
cgeIKghs5ltlImsBS0aJEj/c4UQFRJcr6A/sJWmUbjGhWrTajw5GcIOg52nJGt2B
eenSOZw9OedkWRf+m30JCBK42HhmKBrcUIVW6aZFa+upuoyg0Feub/SznWbPJbl0
LH0cm2PKF5jeCyc51EYDawkJYWQsPllojoOxJyaPUnAEsBOaWiOxJgc0pRS9c7zO
OBb/+pMAzJZVNAmSI76Zr4nmJg1PD3GLHedjrb/HpL56uKZ1nnyuradADaGhvwVT
IC4CSVCqMDEUFe1n1o3y9NjCwFnsymMyPjidxwwf77CFSuNtlHoEPLYUo8HGKjD7
hnBG7N6MyjQkAwYebKSmHKEghcsnQeMRHVbHY7m4gkYMOfI+Alj10KaD7/VXvm0i
0rNqC2HXSpitEe43RiAdvvnW/GXYjAkQC0FUZ1mv9QAUb1MqB3fa9994h4ClC8mS
5rKUhqPtoPyBhUOvas9Lyq7lV10gTnCm0wqMKFxedDooEpbWLhqei6ydoOTCnqZA
RRHoW8ulvK1rwJY2krxgjvm4B0kvuH9lDxGm3O3NllBD0S0C17/xkH2QtyFiSlg0
8aQZbpV1EWszu0IPc+/YIdb+GLwd3biVv6fq7LvVo6nxN/+gTMQTlD7qz+Cj2Lt6
st7z5vuVwAdeMVGhJHORH0XENx8pBNDsuLEWFPEt4m93fgghNic58/F/AW9R6Pev
6Dkv3BfBzh9AqRLe/GEmly8ax7Ebmfo34sFGNFiCD1GuKE2kB5MHBs+/ByFvlZV0
Je2t+zP5IZPRUdVZWEqYURzCR1NMdN6QSbljOvOfvHNuM7jgxbu56WxepUN2iBcZ
A5O8ZQTG8a/mWlpWwK/lYkaQtSbTu3WmEFM2RFZh9ZuWSI6dcMDFszr22jMD0w6R
SKwI5i/6fEnD4zWF1PneFWk9+j8+da2KZFCpIeAYB3ydBhZ2A5StFZzbcxUiSuLc
e4Tm3Re11cVb0qKSfvfCyOnCHxRx2NCnrI25W8VnhNSp+mzu3fnKfNq9ztXZWFKE
jhlO7hLzdo24RTdAr4+qYvukx818+Te81gbKe8yAUPlksSL8BfoYAnFABJoaKgcB
4hGh+1GCqG93ofkAVX32d+m9paHSOjKpuizb8iJcKAE65cXTeGtHcQkqOn/Wunv7
G4+RknaS9CaVMW5i3dh/EnZLxtpjRWbK5z4K6wHoafqBmUqPyRVF7IYktij9Beel
0kcbBtFgdUClTljJXLW5rFZVxVlebAijYDOFyDzqVxUPQizHkNSt58XHQL5d5tCi
LHnPNdnB/f84Cdq2/L1w+3v/lGit6uRvBzwpFyiiqjNNfyVvxo/zkdqNBp0pSfCc
yj5FGjUJlnFvppC6pINn6qhPD98aXZ1cqOjc+yjol4TJq8OEI15+4J4tPkeKWVYm
FERx+tOcoILJ6b/WVGuY9rWlzmsYx0CvsYae/pcXGcHokYXqeIhfTUY6rKjsZ9KX
P4MQjyyJS5Pk0KK6q3+22LfU0r+aZ1BRZY7b0fdO0H770ETERHkByM0SXX4xm1M5
neF+rkVJk5meL+eaCq6+K0wdZ2y64VOzwmrx4VptqETcLKLiMblHigRhZ/KgJUKV
2W6x7Ur7H1s3WawQw5nD+XTzSGn2eds6N5AwaUa7f0ui6616iKB5z5tLGcPFlPjH
c7okPeZ7RfpwopgpqG8hETuQIeMFRH3RL4sw8uvooddBRnBYebaKoyErBv9bbLgK
ihyazRqLUiNEGIhH0frm8uE0HjEZeMinQpFeKcyd4egyhHP9gmEtCkEVrii+zmjP
yYMCa/2kbRv5JW7fDAzqKaZlhBFcln3crlhxSPTAzHjtQIwpuvmmCxjVe0oCoLPi
wYfByxb5M7ID5BTkZy42cpK8cZLhjbLHuTrE7JWK2tWI+F+htzKW5SnJgwECPDNd
YeT4oyA8fXXLjQNdeH7hUMNjnOGjO0QrUoBsRR+Vf2bDFHmDqqaacatSCCGtiSlK
tvi3K3fHigoBmElE18NhrpNZLQ1IwuNAo1kBvuOSpeGsL28PlfhEWbfmaB26yC53
6gwsGgMctTRVBmlxlZ0bXhgySfHgg90tS5a0TCnAlGDkpb75ehXB+Mw5sqzgtWOn
9Fehyo59CWBGg+1p5mn7KWxEUp3hXY3pP1m1aWVEMQIBtTf7RQmsvmsnJB1krek0
TFg7Vvl8nlmqqYFepiw4vECROATZpx/h2sRF7l0Pt80OOtL8SoQB/kjIpWoMFmrW
dlYg/b/me53FSHh2U6WoSDG8aiSv+XB1GvDu+YhfGKyBbxwzsxz4flXdnXqebU3G
KLJWQ7uilczZC/BiAZG5XUQIKv6nntmatZ7t80LgLPpBhYkyPhq4Xrmf9IKGWzmW
SIfkFylhi3wWwDJGckntWhpE1EbUcYYc/cB6jHpUIlb9Qm5W/vkN5fjsWyiajfwl
UXavPf3dtbIxEDmon+VXlcSXDkP6LrLE9njdcqdOkNAAuaPMt8vGdXnI01wJdIiA
qiZDFGwnQUzZJlp6Yrc+m33kcycKOy18VVFl1MODE9cks/DXxLAD0Nja6IpEh3Pg
Qe74pSS5ghcfrglv41e4MEX0OKZVFgB+m3A0pyM+Vo5CjsssMjF22lAb8evZ6slT
DaP7qhkvtfqvV12HgDSUTtrJeDH5DwiEvBYfq4oDUhQ2h1wFlX93eNT/p91vv+Gj
z3WctEPmSpUUD/3Wh1+i3VSSwXbr8cnMDyjY9b3fuf2PqsvKvF/xYDyMWLY09VLp
HEa7Az2lKp6Yerbern7e7P8Cv1PfzAR0iVQjHLVSNPQRSaEdGVAhEgk9Wc48jXWD
77Yz2uJnnmzG3Uf3D3W3qRr6o2eJLHeMN/1LjCKZCf2bG44VsdZOkvlTfVN+ABeZ
7pSn1H2Ovftuxs9NXe2sfzAgNcAP2FHhI3F5JgwA7VTpwadJS/UvDHtNPYCS+0zc
Wni3fKjxR5UuUH+h8ELCMLihxlpLwBUSmimtX9/jmYwGTbyYfW9mRF2rIBQPtg3z
JbHyUcKc1KwfvSJ2PJ7VadJOqJUSw31QZfXSQ4q+Xx987S+v1nVf6tENIUQeb/1/
O1B0j7q7q0fKeqDwmW2eBNihOBt7abHCaZD6cjYeeJVgw+uYkQDqgzhWzbV/+fKz
MUQdNg/YKjZwhdwirNNyOibqSy+sSp8WGG0Yg7ATVJ7a7ub5eBg1sxKnngOqDvKO
k8ft8IApOXLWFixoFPYMSsLfPLyx+vVDL1KcAb94nViVa/2tPRi0gBYshfJCAJ9x
zPfGCOA8bfsxcxzqeHsSo1Bf6Vg9Lx8eJyseCcTY0f9AOfnuitQqw/A2NnCnoEmY
FLrC+iw0gpxJjTpClNRRJrKlz5jYSy4KsMuKbri0Po56TJE+twwqJow4EEy9Lyr5
8/HM0FrOXFBYMk7kym+BrRmLnfLzHkDPyxSk70/UjGjG6gizKju1TsLSIfGL7D/m
X9zqxzNxyT8ZWMZN8MpaDxEEb5vERvq4PgeZpq6jCAM3Hh3QIT0jszDk6V/AmGZc
ou5yn6s+G7VeduTjDl3/nvCQV1YVvU0bqLHMyOTR7BRb0MfPunIJV/61EYGsOuW4
REWdPBMVCJ19ucQ5/lC6TSWSePmxLH0YKI5sNpmoUGczwF/qmhoMLRjQsNDzhwLs
aB9EKPahQDGz0NkHH3XeEXu3IUxTIEtGjTV2+qFDpP0Z4wFr3yX/DOSsQjltzyaP
xdAVo29hwz2CjOS3zLz5ObBz5K4Vj4OjUAa/QiYteenFwrYRY9oTVjsntoZQsgco
m6eQmXIg/xoSameX8ijHgYWnXlm2Irh8e2P82N9o2+sZh7wye0ThrNY6wTKrJm4O
NX8j9opIKf3LYj/F240fuPQbgX10XtcPNvtFwcmPZnZu151TZ6hZxRi/3MXGQbmP
TXynmFpg/MRoYT9/qSnKqXiQLIGpL+tTnV956rVLUXiiY4MpVkftItRebUxr27PL
1rViFVEJo6wNa5dBroEVF0FhL/eclSMoh60UMlpd0z7kFHGu15Pov8pKdkI3B69R
aJdYMqo8SAPa2vEoHjKQeC0ode396K3/bRWsyiSmyLlHNZacGqjTbiF4HcQrHu7u
Va95mDis9kHL3zI2wvWhKbdmrTif1ij6okoZHdxwuADrpUWBtba5aRhc3oZxoJwQ
8C4ZC+P6NRfx4VYUqmJlNRjWd3ZelZ7TjS7LPJuLGMjhqoBMmnRriyR1THyk+6Jn
kTNUSy7zFmHjSID+Wpy0fDJRL0XaBJs8h6vKLvnnIStPZKhLYDert+A6tBUfND1Z
bNaIlwndMx2LkLPnCocm8IH+zKQYUAWyrejI8p1922JNwI+sfwsyGnCyVb15mqS5
pLzVybXCYG7RHl46GdtDgJLmNNsNzuAonptmyRL1V/efjkuu9wVn5wSx9kmFmkyy
QyMnCghM3k3iZKD7xyO1tlz8o2kj8SDPsYD050qZY9gkkUopPO63MTbwP74ZVXhr
jYUnOn1LdrCRgc4I7xCIoboy/atsDq8O9lzcx3PQPb/IgADZRemcIaIg+ZV2msf1
xt92mgez/3cd8CsM179e6xXKR3+QSmDf4tlAF3Q+VNOfkrGmnFbpDjeKd+xpY0K5
BfPvXpxHsYqtI6jmuAHwdMgaJ94q0gpPlPneYh2RZB3bhQedKq6sNzRdR8mj0JSw
s2bno2V+tW/1rktevqoaGb0NWv+33YBBaGny7+UN1ufV92Xbacqwzw+Ynzp7rWgy
oSAUCz1PIZCfqjIec3D864yXE/tCcF+PiKj0ERZ4URuttBCiJ3++HCYgaTcjEc6x
YDRaRsRif9CbwCtxBLECe6bjRAUpbnrAS/aGNso/AIV21XLNCmWXSf33hXwWuZXd
JcIvQFQWTx3LX4pGZjFIMmPS+myHHE/1HdsJQaMeq9W/TyhgoAqrOFFvuA9de4CI
6N0EruBX2VjreGasuuStM0WmmgfXGr28XmUOu7FyyMzBH13S99ipAXllztg5D+yw
NvkxuwdQu8IsXhbVGfOB37IfYeCgjdJs+OSQlTTpkF5c7nUNzJ1GcveYfZcq2JkE
0XKSoJZhSgo3PHuoegR2eH3rRBTIwd/J/zoKpyfK9Dc3VZh7pWVEpxQjDrDpnZNB
s6kM9iztXky0R8EZNALJCHdlQzlJ5xtsL/UaQdU38bJ8TP3H/Fyz6yV9RXNb8elX
gUnfltSLQNttJlpjT7MjhgMpAjvoQAUrp0YGIFPByli7DeJFFAi3dk4N/MemkxO6
RM4Wwp2Nko/2X0vVbLtFdEDWh7RtoEB+6ktgOj9bq5LaiG91M4xt1trWbGu3Uvm+
yZedSfxblLQvs/pIP76uDUa+lrur4gPJwTwVtHtVD89zL9W/d6/B7ppxdWUjq85z
HeBj76eaq5YB2BXUeXGaEXzCux87n5/Ka6JZiNewG7cBST3id2Ms7I1fo80V29bQ
1jhn/Fi2rrmcCPSY1tlWwZEQmq55Sa7jnV9MzZh6aoedOnIBYk7ub71S3LdBZxp8
uXqZFK01/NSrUFUEoquEGQPjh/kq8V3SUnP2DEAgp86sFKJ6hS57BfZrYzUyjQ9n
gIhq39BFInFn6ho3+PKrZAcqcN4O2sxahlKLTXO5/FTJUhsZlDl6h5Gyb3PkkP/Q
oskjNifm58Fnm7oXWlbZ1wI7Fx+plyLqVc9JnlxM/dtiWxuUjEEzTwBVAlscMGbT
Pqn6UiBWS19dOVtm3Mp4MHf08/0o7qxi9BHy2vndH/LZImqdaTOS8ggbjy4ViUSj
Y9/oJ1pn5YOmhjxAV/bAMrx34MKJOeT4Sn65P+BkOln6OOLuP2zDYHmfgn8ZZpxm
zXCs+8+2k43bJKY6c/Rr0YTUnGnrKphuZde4gkTzcs6ZgxBOPNKGJknGvEtVECQ4
mfN71SQ1FkU1mlTGzhK++aDVvE/ezGUc8n0/tnFPVV5jYANTvIeadx0rEOX5JiGC
zV56EuRT21ebWfa5D8pQyzEyCzRK2c7XNAE6RPQG/JMGYgOwkuNs7fJYgftELi+T
2fQ76ZGcUotA9EHUxhot96hqfQOidaoigV/rtWlqZEAD4cph+nBGYkvGivyDnuZx
76503kzJyEyEHEIMOL+aghh+ycPk21U9N6homsi346LGPSMgYwkYoWDMXHDM6KKB
ID+Gb+pQYkLsBgPZKyUU93VsrHa8fiM8sEmQ+3RUBe9OHq4OHwVTf1KlA5p3KaIZ
YDpkjJ9lQAMQ1FYHG83zpaSN5AH4FMz8Tz2g5JMlBs9f2nFVAaulEeXPJBDwEHQo
iA161BDXVOPCrotp+VNw9+xEksSMb1SGn7wz2mP5MspQSZBJDZO2kuCDyiiV0wt5
zdRv41PMgBffjywketpDYgcmTRddTESZ4QPuxAUZuTDBWhizzohXGjXYE69OJGD8
ix2yQULTeIMMTqzz4XXBu20FIRZjT643t/ituzujnTf8B1pMjzGpgf0IVduTBxun
mhizznS+UFkZoOx1yariUPEqlpozG/N5XpqDU9by2VlA198FcUq8ptk3BqlfDGtt
WcExZd7vOTrkYd7jEW7xIUIPQolw7ym4U0/MNUOQcfE6NapHp4m7m+/YSkMtYS2p
q75nHFA64525+ktZTeAj49Y4NHbxRf7QTJYCckRj3DRS8bzBgJ2P26iGCTU3LRYk
jPv+AUD5QNXG1oPin4LexuG1gr3fZV3Oj05NiTtUIsvP11+d1aLShI6fhcpn9uCS
Ej8pEZCilGp5kanK47olp8DDw9Exzdjz66ZZGoiW2KUJtF+zhYyevhRxcVRUkyuA
eA3GvHUrqsnBI92ahbppIdKP6WfQC8IKutOvwys/KSA9059tEhEx6D49uxmKGXP6
oM2xAcL/XkvU5m2sy9LCNyx6lDHnCVjC1wGKORf4erkRDPx97up3CfyDOd/TEWTk
nJI1GGPwdOS6egt+IYHXBYw2iYaNQZyVipRrU968GgYcem8z2/6qcGrP2oZGRwyy
eKuXn0Zc3vr5uIpsm6XKtmgYeBkO7ZjNd9LlycbeoSxYRcDAMamUAtGZkf/mLw+9
BifDPbp8AFHVr7oXOxLvtKZYqMUCPxsW7iAdLzwOdgc5poqMVqRHXFzuKQT8UvOd
RLBe6jhgQdKjO6n5urRZiN6v64IgDn5pzu9Sgl2zLfgGLND4+ELLzUpoBnpAdIBG
YGtKc5ytyR4BfTtMhzy6rQCjIfdrNotPJRtl+RPSvD08NPkXfiEhOQOaLsyBxCNk
0gmbY+UkL0wDWXlgwcsl7pmft9Kw/sO9W/TYzMxgZzVQ8FIEsmj+xXpI/Azc+GaX
tmAzrX0DJav1kfa49pkfQUtBNtld2alBIU9Dt6gqBI6Qopuf892Hmdf6VDl66miP
1PKR0rwVQ7XP1i3yhfRRNGOOBuonY9Rw2+9YwX6dZVuR3wfEPOJDhOh7ecAH/tK4
qwHApMKxjbMxxXz+A+iLaBtxiLfyPOQIwpRAUl8O8pu42oCEp8J07IUHqSm67Pj6
EvMCuVs2bqs8a+501Hie5KIkWarmT03WgQDAujOtP/5GeAgoL82E7hBjzeVoEHQe
b6/HOUTSBvIumtFdBf1QwvwsASAUNN+19XgPI5eb3N/tKcxzpdtJZKxmbdf5WlT3
bnof3i+9M0acwi4EGsoBVxJXzJUvxuAPi8ZZBm9v4ZcrCGbwmieQPIe55c1awIuz
WNBi6C5K4IWKj5efHswtWTQrjdTVgGvKo0E+n9auvTr2QOH/EHK37okAaMKNlI0j
0R8wtrhtDSMq6odxpEzIc/LVUOZcTWw01VeAg2o5wL6to6FN4Z7bQRIBsoA+Me/F
aZ+pWyvcD1wYzzUsOPPdFsL4Na0XE6EFpXirYGS3n7kujD0EiiEUpLPSrcrwAX3A
FjEF5rt7JH1vjQBLYROHtpH1GwjQtKpei+J6CN4tcJ6WrtT/G+xhlYhTT2Bvp8pb
RocGQYgo6vaF5CTl1Tg/8rG0s72f4GU7m6w5NHlkxDqKpT05L4hNduKXhUljYq5W
IDOuUt7PboIVxxlwtdwvboFp4y0ZZXAIip6DEYrcyjL78JN5dttVkvAT1GjjyZ5U
jYdtgmxX0RrWAr6CMUrSOoLBBGoBLXpDpZd+xboue3tSquc4jzLXbGWfJv48mGKV
MTqm7pOj33BXfHZLMB81vdVNhcVMQXRnv1leWtj0QX4ngDc7Uv627fHdP0g8+hX5
7JHuyftL7c/gGTdbtrndGMuXgSabnTKi5/+ZVeLgw9P4Z9l4UVkBFeO78EJjf78W
kO7UQCC/FiFmsgdyZfaXXR2HxX9iluiWThhjuQ58qJPUF/+K7OVmqye9+DUOdy39
5uxL3REOA4zuLLYIllz3034Kvrxrg9/ZjMD4DE4XlsCyB8JTfXV5I3yqj/waD1M2
9r0tNGayiFkz7qWDtMKvNryLQbfoe1VMWVeHkbjPBusdt9/k+O+5+lVE5B0pKg0Y
nuWdIQUso/G8OHaORhJVLRGrMrixVvf9xBkzOmGhDQ745WUedO+dmhnbv4JxA8x5
hXU81Y8mA5+L2HX/V1LJ2n3bkiKyEtr4w6QjfWfCLxuNlbsYYLT4hSqcuagrOBGa
4/q44hhY8hvIQDQa7OJIYtanCNbXlrwZrJ3/psS4Dwv7TFSgRZSfq0z+LU0o4uGt
8d3YrqTCjH7Gpg1NsHi1GOV+sXOP2aUsDcetfGnfFyeGRM7v1rH20H2OYJmE6gRx
BWaqVsih3vOdpJcsTHYdMsOzlDpDRgDSHcDmah1BXmrZibnXg5FCwr+kGR/KsnFF
JSwdLO85iCzdNwfN1T3LAKsXpQE5aTrF5l1PTbLKIFglCCIh3J0mdf2MNYQpzEnE
l5Brqujddj9rt5xgxm+tgFh8qRSX+tG5xn85RoOsk1GzB4sA09B0DxByiluqsCvm
HKftsfGcMpDoHVBj9ZTzT7N8HGAxLAnSy+qaVMCzus30UXVnVU0a6CnM2AheVyIC
V9K2x9XVjY5jtyKboH9rqSvH1mI3zYJXJGBvpo29tiIJp/TskZvMZ+CN8j/NDnB5
Sqw6j2dodaHiwIjpXUPnMcyqmPKYLiLNH6cFprAvlMA+anNgDQ8BtqlCB1r9V5jp
gqqb9y93d7gTkmMXDRRt8MYd5ojExOkZDm/oTztH9dpmjz3yQapIwtKx25TRWLVb
YQ6uAgzveftGrcrTDUMVSDfJ86PrINOttUnracifLOcMgXQ9KrJ4WzajLR5M++vY
0j9ugOwMBs1ouWyDK0iwmaP7b+rZGPCJMn9yRBI0lHUBMG4+vCD8zTtB9kWp1GQw
ykkTPsT3wzA3PemgHYdTxzn5oWQpRwWqadPhNJkZjNuKS2NOnlnZyikIPHInMEgN
ARC/aKM8HzpVQz6EproKAx36Tsj8CDTE/gIHATarjHTCsEimfKAK/odsiUHDqazb
gMNnz8R2ivSbjv2KdiiVHbTm4A3/46C/eoPHn/m4MbsP/Kfrea/6nPw0zWdgx/DM
0EvoVsK4qstw47A0RMkEUYS8EARd5sG50ZqtKd73szoA7dmTqsa+dn51xGX3pGva
HXl4wedaHpaDZ7xLQNL5vUumuJpdek+t0WVLrUsoaqbvwJbM3fGIKCm9T1HbyW/Y
uiC4ZcCFJxUfiOAEB6ZVuN1VGbR4Qd4CcQNR0WGk13v+FFmyEzRIURN7iML6pDKf
mBNH4a+TgtRY1iTzOnRKUFdefcx2SwWcCciZLO1Ib00R9bF06n1R+uh2XB5ND3NF
xB5R25pL3gp1jA6F0PPYhN9J6H31Xp+7WY/VG9I9Um0erXLI9o/PF7CtTrv6zx9G
7EZPWthK9NhjEbVckV8C+zk8rmiGtmoFaIDm32/9len7AhnXsWIG5uC/NvK9O4hh
PfRFKfYUTN5jZbt2RWQl+uKvbW5xgkjWh1vYKBAXa0aAn0vcScLEfRupz/8jaLRE
pyiTd12EYqcAdMLR8cSc3f55rpV6EBMJmHyhDW2jm02ZZTGm7FFHbFdaQaoGfT2I
d+LEVlBVxiZNRZbbvga7s4Psl81tEx9Sy8sS5UDVjJw3Nxi1OYZQhf+JUhBJcxfH
D+92nYpSuOnjKKnPXZfzHnsx/V7p687fNFvEinZSRZcdXU9Y9jGDG9+1Vh3Mv/ce
oBMWneoC5T8EewsGI3bzSCdT3zordGUXmDM4cZh1sKrb6U5Itll0N0MirNeI/gne
AIWriTEY62oSUn4yL1pu/TceFrmA6uF/m9jvIpoBEFwermZyaK13g3630cEECkBy
eK3MrTRJ55+53gult4P8NHTKXtlqAqiU4+W1bbvnbI5fbT3ldI0fWZuQd25+16ID
vATsc3xjREWfkTlltiQDmF5J+YOqP9PT2bHYEq072kL3x4ICpe7u3tGavmQhpVWa
wOl4jpg7zjEisiJjDOlc154DqHghGacim3yL95O1aA7gCQpSZrEVIAnLLl67arOa
LflCQQvwQox9xJmowmbLA6NJ3vt/uCVKKZXITwQYspeX+4XRadxzo6YDBIjewg7v
fjruQzLHk/Zz4gA+C5xL0/WK/f/V18fli15LkfMjQ/zDwOtOZry+xEpCENs+2MZv
2JBE3pnvtTGsLd+TDFGKHHqkmkuYyr6booEcq8p3bHnJKwQtxt0uCc5E1oRV/1Fn
WWdkUnH70nwpGA8vQrGEJhwATZgYTcI9NTnTfw7x9GJPQqut6nhm8nfKtcvyfGEA
Pywvpgy/QdmjJ0QgQexLDQTuWPitiLP4V0JXFWdA4/ta2SYaJq2ybXoVdvgrPuEz
YXJKh6jD9AhmEgn3qWaf1iHku7kDPqsgHLnrj5RT88ysko7+NyU9SvDrdBLEsFmc
O+0U1EzfHa/qDLYlwBhxyaX1oagL00RUtd3b8eWpO79JtJUKLZ94Hp7WW2GI5+LW
75WQXoda6UcHONGO8+aA+A/FXthfJZm10sU6nXcUGHrnZQaXDq5jMq33AmVxj6fw
4bOmtfm0qel1EhuTSJcOHohuJXC7MCqGjPOE7z1e0LxE+dUEuJ8EceICOkq3bOXM
te6aoONjZkC4uP8ecBvv+HdNNsNjWqOyVemurWZZH9wcRIlrsJuw6Fxw0jjkBFDj
fIvRPy5ppDuzNogPVEQCIqfKYRTwDsdmkch+7wwEJD/VXhGO7rBajgri6Z5nFwdM
SUZE9Qqw+nLFidmlKrshyNrzzyjWNIq/gXSsiXlrs4DJC9ejdKoK9Lofxl+CLwhC
Y5NQvMO0+iyj1coMV2Q1EbCwvvTna+wsnBqUvy5j4K31mO/bIePkWfL6loRIFwT1
k7o2bID9KzO+xgI9tM8V8JnWSXndjb1ADX5+JxUPDeKMMq0zj03Bp/NZDChhr0hp
80Eo+0QksSgxlsM1C98W71YerleQ7q0HPRXuse/B23coF5a4fNEIlAC0KBVXhyxW
O9+xxdBCrvLsSuBgE+onTWCnx5EYW5zsRBPhVqWGQvV1Mp8OYdHx6bKXnSBGOaVt
HthN8yj33McVSp1g9GX2ib+5G91cgr3rsc9edQJpZLmrMVp594oQ5DV0bsMU0+7+
buIrYmihdqTB58RLLi6aoNT/eSVRxLCXPElzRYl9XjtAfgMIvMwtirU+pZMQ39YE
ioGTX82lGIl5AkmvLuO5anAcGT6rqzXierS8yhuZrroKAMVnIVH6Ss+Ofhk9YcxE
Qjon/wUBaFSXbaPPbI0QIrNuBh9FvK/uB6NVkEem4qymntxaMHe3HB+6Xm8zU9b2
Ho98fGWEMS/fi4knvQrUv+eagzR0+8kV03XQ+j9bekMWm7ce3lt+87D0QbXoHOGZ
TNvV/erVhW3eKo5j8HKweKIqTlRNhwUoEBtz7imoNulLwqv2ak9LK8AzZZ/tQ3fO
l063spmi+h/KItanxj0pSoWr1+zUqh1eFDDeRA2/6tBbwS7Pq1BRp6UVNaQ99vTF
u/Yge3CwLpzZ1VK8WzAOu5F2ZFp6aiWXfBYCAnhikbau8TZD0MOVXVKjinXyOAeU
CRxU7MsCgIS7ETKFoBAteyqhmhYsTBndkQpL9YxeXhFFO3aXGtGL/hapyo+dHXRi
sYBWPTYC5g5ZYDMFbfVKNjMPWfOm+rBspI2Hajr1IVpv5ZqS50vfc55RugAxiO7F
fl6xwD6txVqImQ2gYNnGizdAMsTtts+hglmDwWq8ZudJ2K41+jk8v91eGNDRHiJN
jUQzar4pDQztqZeGhoDRY7HuMG1DSI91yijCAMv/cshYQuCZioqQKVNYo2HxAZMY
H/Booa7hhhmVvl///BWVB/oAzwZnqMVZ6/pyTDD3wD260uFmUBDXkcl6IqXdkyjK
jjOdgcY7Y9T2O259oJNajzENamcbv5+IuwrB8Hu15vB0bFZKhJcnfOPdp9zVmzNl
43vaSVdDQESvAwOSRW6SCsJU01GFLk+oGvFvCXRybcHM1B97VVoRDHBr82pdb8Gp
UTBpGSAISJPBdki6D/t9Fqw8qWIEzM0TCexSdx5nPOjdrsF0TMzoTvX/FweJH0Kj
aXtJn5SR7gdLY9W9M2rKIw/1tr5iPtbXEPZmrQJcP8IxDsAwiheY8gaEQryUtOwk
Y7gycIzLlr+1d2q4WsLXblGlsLQsMZTWvMSGrN+GGbFlUkALq8zd16WsFNvYBL1W
1ty1Foadzf9Gqa6ibs5EqxqdbXUfgLMhVYaCg85eXaRhaHuf6n99ZT0jBTtVLDm8
0PvgAaPwi0ZSnKaY39IL2NcsEHky56E+oBVHBTw+Gp6CCpLpYsHPH3KhSuyfLnza
wOkPtKHKb8LZd4WEgjCGtW9O+/4Rj5Jd25qrBK2ivhqUjQpHk0hOqL+n4LHx1D2Y
jlufElN1x8xX2BhLJ7kLFCdOT4SoYLffjLidjdxwF3XquPBOeBYLxgtNUB/F4ouC
Q3K0gPFYOhIjrl4/0p/n9FfjxVBefzu/ri7DEF/n4qp6kRR4lCe7qOuIYUUITJTy
FqA/mri2XbRcX1XYoraqyl0psdLpWtcZE9XhHMcOXoOu1t37QvFmXGO8kczgNspW
xrAR3QAysifm65amzawieyPrHEjSiz2IHAAr2qDy9uG5Bb0eV9YDOMwW9CzsOqDT
OqwzCoy4Cwpo0Ot65N3VvIDu267MD7gOVBxtoiuCxQj+DkqQQwdJti7QmqHRBXAU
rha9nJ6VxudxKmJaCOU4mAwJCK1o5qOOgjQJaoRL4e/SIQCSQQhmeLD0as8AG4+F
yl89BHx17i1ZJ30jnbcrHlSw7Kfxdpvv74k02auo7PGIg+svVSoYwRnNWCHmji8c
HnZzDwiK3w5ZDokRJ/KdH6zFHxPCgk+ydq5PWb8zbJisTuX4KjKzY38DIAZ6NWRk
FhqfVpZFevmd0NnCyLgOVyCMzOUPZsJ21l7OGGt7ZmSEVx41ztU9Ei3S64S6gNns
WDbRN2KX/Tk4KxpPIfJogWwP7fhvjoaHPaDyPPZhCXEWjoRrQOsndvG+mtxIC5mF
xFmYPIKIDClgmWmibfBv519Y04/BlT5/n8yEsCKUGKanfzSuitdDQ1Zy9lmoTdXT
ep5WdOV+Pau3SIYpjzaLwMVxisIJ1GuVHYD3nZmrXxXApGiDYWCMQxxi+L9ag9op
cyUz5ooywlpcnlV05RFMHtbhM35wmai1FsmB5kH4uakzlDaPo0+aglASWEGgB1tj
H3lSkevCplDt2DbFw6A+EPrkvVuTnqN+1WQtp8tiuWcqxzCNOScDBfcXiy/UwlKu
6O0FPyl6JgXcNjrGa3tFWLwY5RJzLheIDLMuD0nTX1y03TmVjT9Ga9NYV9SnTo4Q
+qRjNyG88fevar0jRoylb+QElHmf/bYukLrDiLjcg+v4YRa4IU9nu5C4TGDloqvP
tetb9iQAKsLjom6IMMfA/I/52NaltJ59M26vZrq1j8cgkipK7KUr3LdCcHiNJhnR
IHTb5PbsS3L6GahGAXhf6nhNI4ZkiLwYdcWLgvHqZ3eX77IwrEnesXvkdbm7dTgl
aM0JSw7Q1jJ162OVmUT2Dg9ec2dlOKXtWFTh9mwsoFHs1tCjsYIg4eauAKdHQIwq
OKzcenlan0sJfnoZkrmQNxUEimzlMFPbF1R+Sk+XBVa+qdnH+zmJV3M45/SFiwgC
jNsFdokCWhCLqJpM9tLt4uJQRVnifOcY2pBhoEAqGZg88Wt8c4XhChOQVNrV3pfC
cKquWC64vKMfmB+JSwr7LTohwL9mV8u6NcEqKiePPR9KSpipkj1GwPyf8HSRRbuw
3tx3g/H0RP5yRKdOsQO8Ej1QPJmdfNveQbYzHmXAuTop/dSW6CJDIjKb5ww0dwi/
4tWi52YAKwYD1t5BCASR2zed6KqRsm5z2kaMEr05sve5e7g+YWeKhLs48pSIwBh6
4io4L/Cof+Sn3ugnJhRqmhizj2JllJokT82YpjYRzqbR/EzpmgZBexLZEbVqGPPL
IilZZywwOgAdVDGL2MddxxXnKCB7wmAP4dHDau9BFg4jbTfVSsGIAf1GPITkSf0Q
CMdUVUCDt0IHFXmORne6RAeblzvpWri9Bl14Ch5dzW5yKFw+5i9ddncBpZ0By3mH
N7Dfle/MIsRgaZo4D3DrSWi/I1TMCKHfwlmt/sMjKDm33n3Vxvg/ldEJb8aqQVDf
SCi4I+JlYSXJokk2Q2VjSvja2vdOi9KkUVktPxDZGnpPMsY9/CbusKbKObDfPVRG
2FNK3e9wuCHOqp2exmu+0xSQOKUPPA3LU6U99j5Tb+Ntl6B7UTm/PyNszV6oVgkx
Ix3rKOVKyYf0tkPEG/SxyqUXqi8lz79+ZAYkfvKs2N31xH4oMHlsaMH4qyvPxaSq
rf0knHBCxDAvupKERj66FXb6afehf3Ku8Af0k9pjHsYtL/De0Z7L7MmUuistytKW
lxybojyAIsFrZrKN327LAqCmT/EweeH3Xbh/WTlf3ZKQzqSPr8FGGrevS65QW5p0
SZmVyNqmETJ+Svtii2G77vrM9E8zQp0ihEX2H82jq1bhr3LYiupIYmdXNJkm9wJ+
MPv1FIMMxXe8PaZo0JcbRYcDmZbvJ78vkuBkBsADLsqwalCIBWA1bBpi6DB7OsiM
ChUcobkxSIxARF7QqNQnU1wCR0qLqo6OptKcjHttU0nn6P0eiW3H4BlswhFOm/uD
+AZTN/tgHoyjuT1wl/9dIn4SMNUKTVldukEknj7eBw4ueOyb4EjXe+FoEwtzOA9i
8MxYBlxTYYz1gc6Vg2mEBDIMhwrTF2Ooe1COQO6V3lj9G15O58dhYCxm70rQJXeL
dXn/eTS5ZqNXsutAV0PljwYfXxCnxfYENOenN0Bf4CWvJAemvqHcMV6zILrP21Dx
Vn3XqUYozx5JihSel7STxoWtd5nBdvBzlyEWVxgYSau1jTK4iF/mTCsJ58pZg4gO
XM6Qfz/6w1ka9VgXUeF3OxyGEz9v2pB4NCLbxOEH0Xh27UZtAg1jZ/9f8KsMuWXk
mKzn6jwShKKkrB6mPGxGQKUks3DG04SmrA56AZwNnbvSvxTlodnak4wkIQWya+WJ
JdM2xcQp/mpkLhJZwA8k24PuC5BzICsuyT83/viZ/tLUEReanAWIS3P0d4sYA2Hh
jkvM9n+xN9FDBO/GLqPUDFKCYKn4uVnjixS2XteSbm73z8m7+sRt3kHJu1hWUBHz
rgmNNhw+hR66JCcGs8SCnS3klgg8RwNFi1Sn+BRQeCu9jzjUKDJPctY+aJ4MTRvh
4KhyFkih8zzzNVDR9M+V4hqiLVT03QNxRGWIU2GdE7nMhqWJsMkVVzGYNd0lX9vE
mc4ZTxUlBpZ+ve6MJEZcJX6KS+RGXIkbAQpfpAp6xvQYxZSDlGCFr2dDlL/l5nUH
3OcQ55qCsEMb/xJhANNYimhcMGNFaf1ah3nO1uTNzTydQXicWHZ7xtbRUio0uXL6
XcAeeoZ8hHWpK/WwoNyLu/J8QWqQIiH5phb1aC1oYGcBbBIg794iD50Ru08oLQ0G
DBm7pVqXZfwcPhUM3cWORne+acIHsvDK+LKZuz2FbFv20X2CruLdH61sJYyMfMpX
yGsXfo1QEZDlzlXZ8X4g7BXgWN5e5Lvf+G7oIFXbJOXb47QFJRcn3uPJ2BGl+uB7
71QEXFAd1EVLO/gefbkE9cULdMhweKTzt9L7L0Us0O0jQLKqPJb7SedpLxxIbUlD
v7fV5gRQV84pmz18lzDK+6fgcUfRhodpLPqXmtnPrWY7+3HhcMn11r/+mJnUvQOk
jLsWy+hgTa3lvP3SI7HcceDHoKCZv8Z6Z6z2epuMlTxI/LqKgxt10bSY2rfx9/Dc
j7jLYYXcRE223FBNOGUdX/GEba9mDFRdl1t4C2wfPcnFOMDnpRkPuHw4Y4OgZbnn
xm+YUD00GkX0BYsnQl70rL31F149tgNIr0wz0gBwQsRihf2ApC5RHNMxPpm9NMU3
41KaX0Kci1AOjZBOKnRzBrJkwSVAgrIMHs2A8BQK5xv8Q2FvALGIwkFZSLNdDyGJ
zy83rQpEzI4SouuIO/9d+hjObHlhRL8QtDp/4jKMx/tGizMMTHnNIlkkgawmFaxj
I6wuyqNwvquyA1KHAIYE/XvBN65PBAReMCZFlVDYeAHJ0ZTV80i4QE7yF3Ato7Xk
eoO3wuolci0DzqeQ2ZhyZzOTPCE/Ev0cl8VVee8pKo0ZVdyK55ZGbBSOn8FoRX55
KcVEybeatCv+UYA/P+YADirBMw+q68ynGT2UnaNjLdr8OfkGDrSfK6tA2KDElgYz
ODXMO5DeQ5Xs3ZmIQFLRbpgSO/AIIvwOrfzkJIKOI0HV/VCIes1PCFkXCpMf6meQ
5cHhBB6v5a6ZxuQlAMI7Kr+2k9On2CtqujAJjU0hdQoIU5nIGN1GDVsP+FITEdhj
0bGGcy4NJnFYiR9MJUtuN4iiX+t/2yqSfvt5ahQ7EPS2gD1WRXAu0rpddQfEGHzp
QC7O1ytIMdnSQfrV5UZDjaXjRiZNuUiHQa2NKq7MnLeWE5p8F2nhezXSldP5cKJN
dEAi4m/20p/ciuNbbRrP+ix1/+NGIHRlXyZYjPC7qlvYQd+X8II7tOlhXxq2j36A
j8mQ3NVkG+R/0VaSDUZcOQJCXd5UyKLZad2RWu3+YRr3Uh8RKDoRExTxhV/TM9kf
4TTXJCPjvLc+2wwrxAt08vyz5fk69h2rd4KsTRaqqa1O5SrDe/mrTE2rtqTqYVTp
xpV0Kl2v3f4GweRt8k8KW9H/K2T5C4dGyTBzkx2jC0ayDv655hLOgIDsY5ov/Axv
zdh9rosH7waMgN4GGdsINKLYHWDBVTn9t1MLKAzzR/xNKdTxJ47WhX1zX4yehxlt
R1Fdt+gler6Zc43dxCtCLBJO0yrDkdPOuBxjv5j0B82XvCOLdKG1IxbPpMMSU9fE
PEWdnRiaeGlese5+5BgFYNadFlZSjrYqGTfx+HYeZHk2vgNOSJd1OlTa9+Eu508k
lHG30YwZR0JzfzYojC7P/vpIB4ZDSyeW6lMQg5iu8uU/WcQ9MThLwaJeYEtQbPqJ
ttGNjlY66F+dzSC/RX0TJbw01E617gKCkRJHRM2/Fg0vlFFPAs/demr1G5ssykNr
gN0qPnwggqnDrF7d3lWcigKUpKDida8IhTXiwxchy3drCxBouAbkwnD9eG9ChCiW
jO7D1Hfmi8hRjvyIBhz0GDznQ8/nsGJbdUrKfS852Xayh1264RtOFc/5bSAm6cqI
1quXWm2l+tPBsKUU1zRR78EXnx29m+ozKdPJud9ICY17FAKoinqGt2KO9EQnULWA
CUZzEEoIFdLY7ZCrcFKuu38rvsmHt2veysBRcZMfnm0m4QgRIWdB5LolZ02izRPm
QegJqlK08CTfxhroRKcJfXLZpR0BFB4y9PciNfxd4LfmlbyhF9I+UjafEBTHWs//
C1hPW39mNA6UEFc/ttBeW0/A6TrluQTw1STF+FzQeGj/OSlJAOWeQXKgWy+8mWo5
JNhv/GUitK3HtaXq/wh+RfR26ieNeYFwbtiyKaj/LAkKsP5rgzsR5Yt2TkWQRFcW
pArPL0c6sF2VwoQxmHM4nvezyTAl0gQ+r12fwX9b96Y10E8VONR3WTyR0pPGzLq5
lub3lX+L8vlMmMZG3z/SqIl7GJBLqMjwN9yBtG4K5upMzq5DNTWHr9TyvboQXLXR
4iTGyR+7aeIXwftsq8nJDIcyFo9olSWDi7itlNll/fhfIQsP7iAN1WVe0XA0+XwQ
Gr3+I7Z/Ow24HkLzuJgbml/JhHewQFa0TvLMo/6yyEPmCf8Qoq3N0G30veOejTZx
zRzOpQuKy8ai+owAA//l9I8fcquhW+0SyM46XM91QITZtsZwqAvi+Cb19AGp4Hsg
+YUm9GF0eLS557wjbZHXKWsOucPy+XWLViZX3i1yWTJ1/+vNoG9Yxf2rxkLh7ANH
iCfUCoeHmQU0ZpUDBzBWIxNjAhCzpbeu53ai0S9TV/cejFjwWToYyKtBl5l3NMeC
kmP26Fd63QsQGhUihLULw30FMJLLMQqznm/kDIzLNV7HqPVJ9xjA8ytYafBvveo5
1VkQI2FOM4q6vOpF3eMgbRpY8BbqXx1Od4uHqbktV9ys9m9338dhSEp27RBN5x6t
FqQy3rtFT9wu0ZJmcIOlNPyqK405m888L72o3fgTAMaHTYFQZvYmt+63lHUxXyYf
PbBYGfbqzJ+8TSC4w0I4MV9+BkZwHxZHY0ZjB9LRy2dDvLP2j5DQXCtk3fNSxOO3
HH+n9XJybmowLG2AWj2Ack5sPlzlQDS5+cF3p63oh1CIotVwtn7KGRET8pc6n5eb
TyZt3W6zKLE8qqiuy5nabOh+3GZL8/H9edtHqUl85LREdOk6PXfVOyhS9/qOrqGx
QgwSFa1TREpJeuOZKTRi838SlOHBU6ARgQTyPAd5HRRwq4xoWLUoQYKPeDqtXAb+
h1dG0W6gPzIa6cij6+5Ut5VuxUVBM4Cw+9AkF5d8SldkeCj2HF8CpZyL6OoXo8mu
TBAjPSIdjEy4V81ve9jrNUU50Tt/0cnt1KucSJ6o6VqHPziRw0igOi9//5sHzTSZ
9Ca0TLhWCmSPxDYRYM/URMSMsl8HbU2vPsGAowveRm6OhBCItCNBu4yAKkroD1mK
HypzS7ubUPRQ5cSheDc9x0hjiqMbjfV23nb5dpSGH+Dg5IOQ0mSbF9ndQcHKbtwP
outF/ft5IEHyyydFa7T7WG80DwYwh113PWzVsmcjPFr/uTUZ15nxoyc6oPwktUlj
aZMdYxXdD0y8AcMtyReuqtLvxhFQ4OwvJQ0r/BZ++oeiORdMY7uyE1UVwQkzGZuU
ctZKvArQYYrbbzGt5YK4oLZMDHBAB6UXudpcxhjQp4keXIbVO/Phokl21bU6lz93
fNEcZHjosrI/9DLzkIJHJ4gNIwmXWluYLMJ3s2MP7cTf3X4u0Vh52a3YckdEEcAZ
HqNkLy8iaoqd60D2kW1NpbwJQP7J7brKerbotyoIYv8B6I0FXmyCZ6V8vnB6E+NV
fHyeZt6dAPIKm8pZ7YrAHeqr3rA+n6sJBwpCa7pQGKH3P/hC24qHkrC/zlv6FR27
DIunZkw6NMrLP2aa+lkXJbN5tehN1MUlURwqd82i5FbS7rNk99Gb56K/D6y0M9LU
3Gfom53boRXIlKCpzyKdT70uOWAUaDJhurIWW+QOFCjDH7Tsvq++tX2b2DMEklh3
BsbLE4ab/wPkiNBO2JEQxg3iiRJe1m2fy8tS6HYbYlvkPDNXiZqzqidA8YfKw48r
ePj9+zeQlfzr+5lpuwfDD681EIfUJEJ4fWIpZ/rB3dr+5Nt0fBLOkaL7zjEK34SO
MXlNginl6oAeNC/bylWrXH9E/j8U1iFyFfhHxX1O5zIMOo94KidmJ3wORq6lGQU6
ciDL5+i1Siorr7v60GNohUgGrTXE438TnehQln7zX+29HXctRqm8XAKzK/IhDbl/
gUC22mWbs3bLvlMhNYPlIFU++oukWUmREUngAIwXeH5IDUuQa51xEh1LkwU8S8ok
gVyyGKueMdj9XHjEjMhth4tc2KVlO3pRJevG2fBGdURCKpEv6AWNIJMsFhhf2ERE
aDzyoKozbPN6jc5MgNV9sA+NyPhMeolXFHzOIeRe4CkTFAAGTre8i0EDpLeTSQpc
wasr2OGrN3RsBW6NlLLXgM4DVK4W1HBndogRve7hadRqeot+5P3YSytCYv9nY1cv
fWigvgBIzQUpAMv7tThxN3BXmAklD/k8BShs/YL6iLgVUze9RPSqve+h0phslVBs
3nw17o/zpHFbtPDJnF9TCM8e0BmkC4tb43nUe1eGNMa7rIdfJPvB1Eati0QX1mV6
WkG3DKo/4huuzzkywfF7S63pAFHwYJ1IuFC2vvaIyWUaB3kjz1iF3c22doH4d+8e
aXba/WPsjkRpyKrRgNIwJcXtvxiRr6XTHtaW1V6VORScR049QuKROBppgifLgoTw
o7/QYdl3+AQAQNuJSFzCmPQKdO1yO/QFpLFJUdOL434qlJ1/FFOCZi1Pv6jznuHU
8g2EZ0SmOoUhbCLRcQI3k0M8sDYNVp20N4zNuW5den4RoCgSQFdBO2k3bNEsrTnd
LUpt07MB0Dl105Y1O+kud0ntPEe4XLlO2pt3sqh8PKG4one09yH0toidfXCmyq1j
QF2yWHvzCJdTzDIFbCvIfuX0c3fGXftaOUeHDlL5Mxv7V9lPJNUHezj1nispKxF/
ul+SU3FYMTA5qw4Xq7LQGerb+N3whg9Tek0/bSn8XKgemINZjbPqee5SmWYEcxa9
KqgjJbVJe/8JKVYWwuvtKmLmEARbVJulXwAi+NMdywS0ptjMB3yxbOaJGCZm7GSo
FHwfmiWofNbz0nOSJkrnLobTeSkcGgk11+QgahE2WhaH+LYzD86oX3fIFeJJSx5/
Mq+at0L2dOI0UXHY/i6/FlOsaRa4Gv1i8uzdFIB3OMtacMQJ2qDperbPju+GGQ9i
VrBILDNHHlKeinqyqDYnOqyk8zo3FCNY0kDBP75PMaeNseeLdqipham+78SPQlaT
99CSa650XQEUJiXRlPQn90VM2EiW+hGM0qX+yqnlP4rXSI0tXOdUx3rLGV1wExOA
7G71rTuziLMo1v/QIfEny6+MOQMLKw5v7M5AHapz0zw6Ap3gGZoIHqNMF970MsuE
xa2it9Yu1/oNmrTqtG78PymC4r5fVZ6bDfjVC6Wj6mhOCV9EjAKBuD6H9c0xxGhf
IX0zqRlx8QkMwaxpLzo1Rg9VewwYg2a3xLZaMvfvp6QINBCcK29OT0J/kMR/dqND
Cx9ac4Lty+mzzwVV3VYhjmWS5Tv/ffLLftyZQKkjU9GkggARndsZsK41Lqe2cNZh
IcVjVjeaF6t3vn5jAFphAdPUt2SBvsDitl3VuOX0CewVJeAG2EFL9UjVpR2K9izc
mRtYc8e/QMWlALn7m7wib+l/BqM1bD/KcUicOMsntg+bigMH4OY1HOKwPz/UrLfT
WKFCEsFvy/ONvM7cr8V3W/miQfIJlZFsFIgozGAmhBvYITSZNMeqQV1Es+Ib3PdK
S4v5dW224fEDY1Oex8SxWP5COZ+rMPRB7JAQpwVkJg7N3jbDSUDdTZnmf9uhP5cN
JtvaMZspm84NGTxJ4dm+yBn8gejXX9UwFkdzz+QrL3ynrxJlVCqh6Sf9EG4wdbwC
/IQA3GVWaCiBJleWHwR4eo6o1dYNt/yNWhJPPyLYnDnUaUB7rXR/VBcYoeDS8aq2
RWFar+swwePddptKB7ijCaSr1o3RyLIXWkXPcfd/hHdC9g6QIiKz24OUmwHg2MhM
Sl626XiaYCd9b4FCdCtkD5bGEDQ1sfqwQejAStqSuT7XEnw6aFGWmwA4ikzX3piT
bZs6FyYTg7ss3KizB8Bdyxm6tM2n2foolg+cGBe2SoURyKseIiARO0m3W2d4yD76
3w499H/gN0mPv9FjF9kbp2VBfMDh3uaxPq5CFNNyGBuRninQis50JRcf0Mv8mNeH
fRg12xLyekElpFWuRkICllTzEr0sMC8oYTMxSYkuEmO+cSJSS+e5xcDieBa9kbAv
n52j3rPjET8SZMWe3S1tVtn+ZHWwfL7qzJlm3FeIL76TMGj4VpzATDbm1ROvM/gJ
LFvcR2t1dVAcqm3iD4A+txYbP6uzkYca9alKGhfUu0qUuwTD74fgD3Qhjc8LbARk
CWuzoG1kg6mEKW2PRPStRek76Kh77iJv4fQqA9FETJMCWnBtYGxFlEKDblnDICbF
czI0jQz2Fvsu5FIIqG1Bma9eU58p/n3fb6hbjJExFUlhe/VH/osHPhoCseXYdbWx
moCkdNLHVZaOPHZRNmVMqe8MCuXIv1Y6we1l2q0KH+IKyjlvYThSsyU8esMgmX5C
SQn6VwwTDwxyBJCzHK1yEm0SSMkM5A4TmLFNoraZkiNROtZQr12y8r13e93wsx8d
7OzNLrEa5aaCmQ2JrWWPnUXvJJIBzVwKSiq4rx4bx0MxEkLct5Q8uH9veJXkYwM+
JX+WKTLobPrRlGTSAFeldFvkKp+wuNyRpSuCav27CrG6UtR7B37k9ZhQ+YBznghw
CTCvdqD57uYFtuoTklE+9O1c0dm+9lS7C3UR2HdtmAcox7TG3mX3UFX4N275L5ul
ibvC2zJvsbeAnbcx89zFrv9VRz7qF2lZYzaTp1couGawyU8SdQH+NPGkAbWKm1Ex
2Ma/rtV4CJeZ+g9f31Yg0L3ZPorQxpFd734sNQVTCndaeY77bvM+/ItDlQtyaoGH
bee6Zi78pg6SWENfYSYs13feHTaD70cKsGpjIB3bLsN0oVooFRSdlUVd6+1DprWU
RYjTRbWrekGJMFM9UWMSCQEQnxHeUzyrDwST06gavKD6h9SvQoRpN9sQOdG94Pj5
bKqe6nxgzoNtGET0o6bJa6/0bJ+ID7yoo7kbFT9y0SFwlAtb+p7PUrvRZpWWNz7V
kXwm4PEJYVRwdT2Kq1v6bSTbIXrijJGnAlTqCgilenEUS35Kmq0m6xdcNxSMIKoG
bEhzTYObt09Lyx+TKJL0eB2ixxbVWU7Conyt0sGCesMudiJt90l/KRuyNqTBUfKe
oo6CEdHGMZnT3zjSC2Dl8BP1CD5o1HIFSMzONuoSzlPC9lFxq3eKGmItSAw7dtho
Sox0ZP+s5XudB9s8oGgkpxmiCTmUVcbIeO7SX0o9O1jiHVtVCAG6X9PK2alDRNsY
lIAiiMbus0KfD853WkQrZR/Cv9Z2nnjeBaY9CsSoAaImYzs0NVz5caIZd5udV5YH
TMmbHbcNw5SCZRENK+tVVZict4/rNQrV2ytvXvGawbRwlo19lObRYUbmXtwvJtZL
W2bA1qs49kB7Rc22lZ9Tr4AD+gNi9BJOTK3tzI98Ud652CtQ5F6DN2fnlibpa0we
XzZrzOtUlErENwxgPphjCbMvsTfKwgHrXaR4tjWKAXSAvC5DmfAxWQe6viBxa0i9
e9JQl8bbyRjqixw72WWeK4eTvK3gzRUVbBfGW3G2YmK+2UTbv7FghdCGvQTHKF01
j+0Ep8xp1n+/an7fxf1V4zu5sVD2G3OH6DI6GIYELN/ZB18liXacwl2kcrOwVBgU
e5vaHgYSbNCs8ffaYShfAISleweSxITjaD2cGywvotewmf/a8UgO4sPdWtd0AjLA
KUMnJ+9f7nX/9pNvi+brsCBmPu3z3Z2XzVQA5aCH77DRV8APy/JaGPwWb+DHW6qT
ARTEEYm/5VPi4BgJQPmn5E6gp51U7ytGb2xTEM5kd4zt8UDRvMr4I9glgqVM35f1
QC1vNGjmxpzP9UQm7LE1oqibGmNcoMGIhSay0zZ4MwiLwQe8EwwXMrCAchFpGPkt
Rrj+91U7awbmwXDXS6D+DnbVEVF2Q7L326woyninF8kK6WMLU70dF3Scc/0te4XU
FLgcNt24RwjzdqWlhPt3hESal+oY+0BHQZlhsmCCtg9nF7g8hC/TKzaXs2xPt6wo
5ZLRW33NFLW248Gy+WbjHC6NYGtRZcZmw8fZraSo5Wm4CoXpV0gtWT7GlYDFObnk
ld4T7nxwInPMStSWmbvgBXFp/l0td3BV4CtdJcIt2sJhVW5Re9i1p0H/Ogqm+AMV
E+oZ2/PTVBF+Uv10SvNznN5FMdrJ+iUgCbSFb+z6PEqrgjSFTwm5v9exYEy0BHsC
HQMUVqqw8DaUMoUmrCQIqx8HTsR/rI8EUpMQrmQHYQGEihod4pRTEh7DMyyoIN3Z
jGOnlTbutv5ZyVKo1YXWhyRsOCjzcz6UebxndUs9LdI0RQuzxxBKeG1eBxxvV0Hp
pqKsmCJ6AV9RxkIJX3OW3aUOCpt3iihBfSt9stsBlMjmNTgckJ3HpxqJ5ZR3fGou
0Dzyjr6xZVbMnvB7yS5A+Oj1TfOgp/+7RQ5X2TlxR5Kdi5076atl/3kvEsPTy6WF
4n27dE9qzkoO7nM6HPSfeNNP48O++qwuRA+ggutOriVQtgMKxp3Fb4L9yM7mUihF
TzAzaqONpCKUXBLPQUyPUiD9cOewLR4fIwlWsqWwJcP6XZGe4Zc/aGcrHFBW0Ixa
OBrYhOIvDFnMFMV5WQOpE9Hd3mwCHOxUuAMJopWM3UUfDbfacKcziDyaP7VB/Fc4
+DZRsrg7uw0vXwKKJ+yXG0jkSi7TtEnrurRhDiytOqADPtF6wNTnmavKPZuOZzGY
8PL+q2BVbIQ0Go+xGLAbOgST4rEgxR8UDCu5xBrH83FIt0I2ZEcylayuTA1Rzq+7
IS28N3wBbOw8fmGgw/cLoZLJaBDs6FjSZD4kre4y5RVnV13NiEp5TbDTUyLfzTeH
9stGuzSbEr5dh/QCv2teIQdAe3YSqAYD5bAgQAt9wLQ+eB/N7zSBcNsdvKZFdexA
/8F7sUc8HTwaGbIoUFZdKY7/4DxIvRI/DaEOKKtC+5nmKIFM/FW07OW8Itfo80Q6
ejqL3tSBwyb1EOuYwDCcyTKHOFL/GXo6EZYhqpGU+KIRHqvASC1OZM7Ii1qNNTop
7st4nnw3IOziV/h/RdDUx9t4Bhvip2uH8Dg2Q05uihkb04juj8F/fcPqdeB3o+Be
Vg0BdMlLvycBH2UdD46jOTdnrRV3wJ6aErZcjQzA35O5/BOpexeMB1ZpA205crYK
iY6Mb0nMLH1mrZIwzi8nbopL/9gI7hD07TjL0J2xer2WkDPyhuQFdoAOqf+3LlMW
KIzm8lxxIYGtktG2S5NLb18ZDS2NkBC+VVcS9SxdtocyK1E8EcD0Ki9wqOkiPfFG
Bjix81TTZRfZT6I8q7j6aFmYMcs37bqIyD36UNAmH0gGec74LmqlNVS0Gciis0oE
uwNZxQuTkFxWTKRokc9+wkXXqLOXYfmIyAhVV5O1uFmyMPAE3XdpBfNRou1ctNvW
d6y/6hhi6RJCJe2sMZsi29MHhqDZDmiIda+akliYGPlRSL1p5VH9+JCxEcGyvSDL
Ro3XHsquaavESZctj+Iup7Gwk57Lck482Sc45VZ1Q6tdzZW1eklhl1y/6XnVGIgc
I109oqZPQ29t6aluKtQITRIwck9x5yiRvsb84VKHIdcqqMn6cdmUH6eUvHwmLdmh
VBONoP18G4OWvkeTLL8cPZYA88+5FYaKAgeK9gd8xJAsjvIA7Fd/5ZnCgM6yIRcv
yZjHbOWmVKsFBDMTL10vEad1PiNN4+wnO3ash1lPOFGv4Ib8D/BoEvshvc95KzST
tt1xvJa31olOf2eE8vJuM17o5mDG2GLGRhE4mJuQqQAUSfBdJ98vwSi4wu8KJoXt
OE7ZcNVpBcVQAJxxmWCJojJfZM+a+nZ4WGeIYQagMCCMhOjv6afHng8+oay5Yszk
i6ysuQER1hwJSrJntkD/OcOWOKtVss6QaeXedD1h7KQXZ4onRsLbZIDfBEgACMYt
r5Zbxj6tfvjYbEn+3lV/GiwBqwhVScMu+KlOWqfuLXPUou4a3HitSAmXLn+vds6G
giVST3hSFm9YyVm8WNcnbqjkLHkbl8QNlFXV/2msqLDwXxEsTjT8h5MmkiAqz0dm
7Pgr5ZJhy3gMETiibCDwn95ZaQVCXDRBVfxwRhaPXyuJuAjNdTMns1GcEdwZt8Q5
f0ddc/ntpe0V/6cU0mx7OXcrui77lRfpLYXoLSKJW8hn9BcpVpZRQmJx5AjcQoD0
Vyp3K8mIP52EL0cudfpvN5tjjGu+Rgt3EFqDLNzyQBZD80tS6VbH2F1JVrnUx961
5Qs8RhlDwwFr879dJuyVLTsyz6YXa0qEiccSO6ENtzX0bhW9eoYRZYik54xdj5sa
K5hDC5xBdG5TwSC6qLHKbzwPhqi37+oGouJuG4mzhCNCePmvJtxTSAiZS/feRd6N
ISgaHuqQRGNDQc/exoUITVUhMkV+3gN3pum+cWdJDPKwJ+f3USoVwlb+9Vjs0gzL
PdRev2b/ExVRYZToMKHrDvEFCw7bOOJ5b/2BhtcuA/+TpDF4tsiM7tlqTwmxp9Et
DD9AOmNw+pUlc1GazHCI0JZ9gqiRY1oky4RDmZ0ZZ46cveaws7PPSMzO6Oulo0RN
5R09z7LBKhAman+ozH5JAmbQiN65q3G6gqTpT5rTxKJ5QArh9KEhhPtGy1NBg26j
vGZ1MHEu/FXXwVj3USofrnRZWCN8uifY5xgEGVPdzGEFNiX8GOz1khVKaKUb5pCa
aqUvn1+UjzTr/267ioCvhrnro7WiSEChJi1R0OS5xf9VM2DBCTW7l32Wv9oXeXyi
chzgcYyPKEHwmcTsQvGgMLx90EpXzA+pUVIm43R2dhFZq6w5UJ8S/pwrv9MjQ+GN
zbOrbsWHiFglUwe9skwnZ0rsbJzXX9QJSJ4ueCFglkXvCbzI6iMmt5hH4Pn+ubru
REXXfkAza8NJRddfSXzzqqwIu2nHVM/v2BswXff01fgp3VVyUInY54+jWFT0z8Xl
T6JjfDvF5e7f6pglWWBXUURmMTYllvXiszUlT9ybCEMGtqhuoAlj4jzMPAUqtkDf
xAtUkFFu8Ajz7fn2db9zbCsUj1GY6SN8YJnXFSF5QJ2cRCGwM+M7NoZNREyZvEC/
MlDHm+SCtqD90N+7S3i3uB5Ezqcw7nS64X3dC+K1MN/LYh3VY81UGIL4H6fuSlxm
UptZ6yUq5RgM/oMIs/3Srbet+mGs48qWUMkUEMWv323pn2BP4kUrstyCU/ae1C5o
NJrH3tRyhLUa9sSnDgFzHYgKsCVerCQQwVuF2CxH9tNs/yQTY6Y+NPt8TWfp/TfE
v2YWLPw9XAS+tF56EUGB9dhmiqJcUd44VeXQDeVE3IefrTxDuCsMtbo/tf51hlhq
hOVFm/VW/xgqNhgaPfrp3YKeGnoObjGGakxrPCmIr/Vf6wvEJxIjMvhxI/T5T8Z+
Fnlsg8KyoStgS+PohmLKtZ2ioFSdsHr/kz3JFzkW05cJk/Z6o2x13GtHvC7aS5+2
mVQW358iPN2h5oXgdAFOyhoPQU+c/YJS6re5xoa18NPNe8BkWhNzBtrgEoy1eWRO
jY5cQ8xxxpg+SssMWymEAAjbE5Xg2g3WRzV+Peg5rKm6M+D8pObLMeKhCfueAAph
jzes4zq71mKyKSqDtbRPBZ5offArWRXcXOltjAeW0uMltRTTQNzh8p0G97aoXyvc
xjvKHihLEtTQn9IqVfCTQxKaiHBacU68rNd8O3hWNkyX+V1/HukIz7PLNCDsGHjf
zWcNcAhI6MOIioBzs2plEVdwn2Gh0rQoN9K+I5YyZbSj73nKzESzKsX28KAha1lJ
1ehZ3zyz1QX6xv8a9dhUyrPBeFNviG+MC5ooh8s18qBl66ru7jREbJz19zuGGVFs
79NIGtzhtjK3f+KOLMh3PYc3BJNPouHhPQS4qwWET1D25X+L0ryefvjXPV7tBQG6
4J9AnjCSVIT7hojXsR7yK3bJ7DV+vQjitgxBPA4DjQ6Nttb7m7sdPPtZCrQ5E0+T
fAylMdwWtGOY0LwKi7lhAM8JVhwrFagfREOb/ThsIa/GEhzUIg2VLOjsMXwvGdmX
POQHwPtdxlyP5k3U9vf/hCi3YbNCC1tm9eowgICOOGTonYzHEWv2P9g03YwQvdis
72Lb8q0v+kLm6mqTmo3kLwMDw3IdaDFfZTms4PbtJOisA7/UCrB8c0NZ1FNKv3Sg
PjuLMKTcE54Llkniwlyp797QdzHyDgUw/YUz2TlwOzfWlhyxh/opuxBv7B15Swal
hddWKvgj5eIL59fCHdrWupU8AwL1gOtEEShZTGHcmiARXK2gy3X0hA15cryk+Dje
7anr7ru1RGys9FKC7MRA+xAUtR1TQ4gBvgw59KDnxssUSnCNl2r3sNqgSH/hKc0Q
semQpOJTlz/kRGIug122QKGuY5OLEIm6euZ9DvPrrw9ev55ekqrmTyNeApjSrsaU
fi6NmsBsR6ed377yIyGMMA1/uyfTnxo3jX9+8tlLMkicMtgYqV7lFWmQfpio0tBu
3Mda7rPKhDoH39xHwRfrPn/zTkXhll5yAjrXqkgC4adprYyvbctEuF2SxJHORzCg
As/HcvjRwNCprlbFiJHjcURUAZ1fHckxBAgCB6qT5pApCNVZuhClz4KNCNnkspWM
jZxTUIeC+GGsFqIqJVEy4fYAe7ek/ZVy7wX3ig+JOHQdb8rR+ePKkO4fYQCwDQCM
epQ7uRJQwDCAcNRlr3EJEhuSq8GcQ5THr+roqmd9WSAyoj74HEtVkkBUGCRayjOa
T6H7HYfXuf5Fz2utqiLU+Lj9LwfmLWWAnt0/FgLUoQUk4Lkkhqf8M3Zw5jgO7H0t
6+rcBRhI8zhrJXP+1LG/MJ+vw6Xl0gKiEQeQkJbyI6uvjSeG5lMh4E2MQYscWwP8
fLC7p26TG5EZShUDWEb82Mzkx3iMLVyH0gsbxitd+NFwIfZ9HKXkof8ZyN5ZAJCG
4w+6EaGkfBDPuY9+30x3bjOC45bxlFujSh/wHMmlzXUqhr/e8jaoIZYRh1rAZmEU
IA9lIKurqNLwpFI77RhBptOrmf9Pps8ATNxAEXqKFZI65RhpInp97fsmZQSHmArE
1zP6G6x/oplcsKYw6qatv/lovQ+2uQI9WVvR9Iqspf7nhwYY8/YfErXLgL6TbcuA
lnrMLRplAEdN85c3Sjjt6R3JAy4DgxJbG8sgGRflyRbrn7dNERXa28FWvNzDOwFt
tdyt8wVUvwakvyOWU73VTIHBu8ck/OmLmkLkNb9AfNE5VdeahWaSmKlbqjVd8AJZ
rn1igcDYwG+2mFVsEKhqoaL7UxzOvQ2GgT1R2s6MGqAIvpLPrXOjLSe3zI5RYyYL
0VSNksGihPkYxbIgL6tkpwEJx9GoRMgGgdd/M/js91a7QbfcM49MnAXUZTSRtmBP
hJDYA+nKVSYJQKZIuS2LN2MCxaFXWuxZnZx6wie/adRsZ66i/gigBCzLfl/6NhyN
4TiOauarHuC9P3KH8AL8e5+sGSC9F8SexNMAvWikjWS9dUytDxmbHdnRgioO/ajB
JQUjndAvx3gnHVX0uIPrvCO/Z3FKVODSsTPYzpxG3Z9knmnauH3SqXvwV8bgYusI
UBneGjX2fal01cNM94uu66BBUiTq6YrFUn3pIoNADA/gLDeer8ttuM3WJ2g3Ozzx
8DeIGeRNDzYmCmKERBnB+cX65qLUHq7WA4IJF+F38tBXgBXo425ipm0SZx8sipPu
RDxlvyeUjyqvTTA2j/uRmIwcg9skMkL6seG515WZgGhkhMbqjSgEZ+6EOZox2vmr
qqV8Ynrv4ALnkIYy5Wih9PHvWKHw/B9oMc4pWx+X4SjtMKJfP/vRcIWhxlnx71k3
wK3SscZMttGCwo4NxC6jY9CTyTiGRgvY+QoyIrWFqifaU9eguTS8ZYeBO0UpAObU
QWhm3dJIfPpareuLssO36U0PFCbj0KQjnoSp419cYA1GzxYudrdu0Mxb2Z4cG4/1
+LF0NdaJQTVC+sHhjkLL8fQjq82U+WaSdcClFQC03l6cDaZgjLd0Hz9v2U00VKp/
BoB5hHVHHJ7UcLxLbdtR3MNISmhLho/uEY7zd7DGH0OAwzCbnTKkqEsemtOsLyjf
Ntxsi4xrB3Gkh0VzMQhRpuTYrNU3PlY0ujvrKCMnvqjkmq8xNuaIgFdArTXKl8Gg
5JjkMBn6H/UzpYih5YlwWr1D1tlCYCh07+e4bLB+VaFuymoFwgKtwzDbPXzXL6Mv
Aiohtw/2HKi36q/a5/5b5MYchU+iiSG5H211xuLpHicnXWn8NJCPdnja+2nb/HIf
uWYyn/HcHFFmycF4/jVQUb/Zj1CwhH/e85AJ7RxpW7QsjPDmm5vsP/gBR1x+f6Tg
klW6/Pn3QwjFpPK+u0CfS1wKLagPK/rgMkljO0jSustN1Uc/W2ckF40KExkw+khc
HVsyLXFJftbzHIMLJOXYYBUXCazQ2AullkPZpphUD+/PivoIIZRKc78BhMZF9Nhc
1h5Fik+gEDWgGE5yXevQY/O7MffdxwlDbIT4Fjb22REmARzs/6lK/T2ICzH/dYVy
lkSgmFESf+awxRZG9bTdBNYkOExJCaH4UwhIWKu3YU+ozbO2OO0231ozvg2s0zvm
xnEpswbvgaIUZZpIjPhuDM5eWqSM1vASi/gsABW+bpCZQp7GhMwHBv1OLTBoQ115
EMB5YL04glyXP0lKCN3FkxhQbTIAu1RDUPEACVXmsQpOzw2hF76Di/ZLAb5UE+Dx
fKYzE0A3Si5NhzGJKOUaqUcMbfyIf79aIqenBJ2akyi9yt0oQFGnsyH7Gfr+Gj00
qCZvoxI3sei8g7lqH76K6mjEC7k249h5t7XG78NyTBLJ9mhqa2yqTkLTW1Rue1Qq
T1hCsiTdwbuj0oa4N6Bpq9Bi/hRQ5ETeedsrpLwQJ6nSby6lZDn6ECW/thmV27x2
K1PlTmIx8bcjo/IYUJQmjFIemI7jztqqy04/a8COzXjkgbywNRMk+su9U7XswQ5w
WmD4XNR0ED+8CdRmQ3mzE65LQDHpGOEGWc+NSdDfEza3NOFRcoGHnRQAGkJcrDKl
d25MkUipv9sr8JfbkImzKVDo4RKPv6f+4mMqQiV5B8wK9R35iaSWTFjHLrpln/UG
L5TEvr27jQc7awghXvzpo9/Jo+O4q6245hRGkb/LMPfnpck1LyXyik+w5ecUxlnw
uJyudoUN/WWo6bIij1GiMAqDH7kbyhNm2zxlT+Ud5xOZ/1w9i3D6e80RbO0f67qr
IBlDQ66xTNtU+hKFQj0ySVTFbE2I/2Fhfh4UnksU/Vp+Yvl7+hNcGhwmoprv8JG5
aWEzx4osVGpXVeTCBV6i/V4lyRA/bUFHxXUCFI8yrADeTsZHJ144X1MBjWgMukjA
iO8ldvqIAhIMRFHDGAMwmXS9jFBkdRJPmuplT+vNOmB+TA1RKAufyJG7KCmKPTPW
6K5EK3MN/LH+55aMuPqUZiGkec/BoF6vhGeHMAcFdypkTvs0He/7D8Os8CLPHqkU
T2SRX4Y0ilnmQA/t0ZSwCULYfNRCJd+wgylWuEwjpkftH0c8NDkNfgpgB1hmbYsH
RyIpOK2nkEdeueyMGt12+HRHg6YYbKdHZXwreVHMgAOCohq0Ly9TC2CvWAqcZUXt
c7+vkfXtg8RePRjsOAFLQbvczggKBbFVRGYBkXD4bO5JSAbFtAlMYLMkLL+mlGHD
DxguXVByS9UhMZ2xbSO8YH9ceZQKoUKmoTtmueF8r4z33MZrKQbwvKqWq5QuqTuz
Gpb+bkVHwIUCiqljbDvV6u7pomrGxiRCXzBvozgNokhoEJ/JWaD1Jz7Q35EN/v8z
H6NT8/tLjJIAG8ZdxoAnB51yywfALVzsPXCl1FULoiyzotNMUF5e66U/P4WWcxH1
Ncsr6noLYbdWphEtPPih4EM3atBBa7EMkZIrMll5bec8xsATBU3nPu5yM8Njc9q1
8E7W+IDzdAOhkCZ6GT5bAf7E+5+YojfBqVOa+bGI903v09UTNZXLlqTS26Ii+ys4
DKpu6Tbij4A80Ct0Jm0N8P+lq3XtgmXFUR75TcirOkDHH0EtaYMQyz9HilrpC9VR
9HZwoNdcHLg6hBa+bHhlY7mpc+xIXnm9Cfp06hVRgjyr8I2Z+nu2s1YD4QcefAMT
5m/0yJA/q4unL/92PTeZT1xkkgZM7TFF88qzilInZ4UCrBy5KsIV4gL1ks0pVoQT
8gMHh5jSjok6HXyy0vhnj7w8LBRoMrqE9vdJY2ljqr6IymtU+FOJMfSm5w7W4eqa
fUxdwEOLn0izsYqjo62pHdamQMJ4Akr5W9tGAyBgpS5Ol52AvSoxN00UByclyHTr
lV7SV5wqDdeVF8vg1pgbXldMsCc26t4ZeP0WUBCcub7D+qk/PrvQUlYzs7YaUAiF
X5zEbdEi2KalLMxoBTYVPxxr3fh21a+20kczi/UAWT4Pn8d6Y/a/C44V0kIbezt+
W+yM62qjWQEfIYw3/6v/YJcDlKX6eEze4S4qU5yEfJjE3vx0vEYXvtpYJ8B7urvt
SoN8LB4DBWLJnaykDG2OYpMM9GmfRHVSc5MjKfPIAtYdsw4JiGV5xXTc7r9gn62b
RUfy3/nqt+ToSlO3n0dE/xbdK/md23XvG1SB3koIQsZaBC9bdhfqCe4o0uIHr0+U
CY6QFPPBAEzbavXK1f9jc2bK2HAsUjqeMJEgvhSIyPNRZ4qrUda1i1e+iOnvb9Ug
r/+ZSpAvY6tsqOltFa+fyQzq4hM0lfvxM1P9WSMR64LjtYY/74D5gNi2b3MfCsu6
CHephrnMrK6DLr5kJJCyvWw2DGm3Wxl/ml732YIZhNNiM+MHj4H4wazWPy7VP/9N
uIx0a8Vi4tQ69ffnp9U7jciB9+Etsfkt/IcYD2rwyVJX+GuoZSb7apSHDcbFPqJq
fAcOzZJ7mIDXFpphx/mvKvxZemvDnqsDTLtfpFDGcW7wPNRDJAlo2a26vuPPFwwZ
GVXHpzYPg2kdkkjij+OGbOWmswjAWU+SVRIrrUrMVtSx7qAiNow7cbDEb9r9IHc8
xyzhBXAxf4ngh/A2g6DXo2fq0WJFqZXbqYm/4D8RVYvpvE3SAJz9/jBUGX5cqh2C
TVvbuNkUiCvg9L6N4rQEP5MurIiAT2uhxWYQKMYi9JXBqt4V9nDW2ZGPj7GjZ5Xw
48Lvzg0HENZIBBdA3apdx0h1kAjpLa/ODN1/fkM7FaYA7hwoFwrFqXvgneiIdgwU
klQjvO+jYuKCrU+0jZgvN+kfpy3pdec9ELvpuMsV49BAL+/R9FKJ02OJEEi46olh
44d1/p9GgdV4nxGbefbdUbk9v3FUPqS9a1qKYnFXv2vgOjKwN+WM90xwlhsnDiWa
lMruPuhmmFQTJhIfuNQmHBiUBRly0MB0CbapotmzE+KyEPiFU75d70hHc+OyC3K2
jkZE8t3Vy7y7N+U+4w7MnEIp/zHSaYsAzpAbF/OFwIqd6QiR9XGAVugFbwb1qwgT
gRuOFNrhncH32hB42fIPrqyCwETpuUBk4rnA49Wf7erJelrC0SjWhUIljR3GOMhe
wIEitD7q6rFl1r6I9d3v44Hb4/6lo7qyT7OqBAZ7uoq7M7xmC+Z9wGUYlWBSSqCV
dtOviX2/TuVJ+MwC3m5XasE+twrm7nH8zY+NdcajA/c/ZmHq+iXvlks9+45sjj9e
XbJRYRxmgZrFKHX2vh95Cgc/CZj8KCOsYMIhdZ0hOImhglwF2adygxdW1regnvXP
/Fm5aKDRNQtv50k0RSxRN2IjlVAra/l9DZR9/zRGH3nyAUglsmzTHHSZxcxiS3Q7
RrlYmT3yfwZ8XGQorIazF0vSlAoWlzK8vkmpxV4mDipWOJhmolBZWYyjDi+RInWI
gK/NPsLRX5Q3k1jl2XNaUJ4HZdQh/fjY0MeWlS6gzOAEp2IazIJ/6bAsIYibwNU0
YCrEylMTJgo2pGgILZMsnq+2AXpGHTdx/lnnorbNxzj8nLALXqNL2ByywiGAnTqO
kkP5Fj567Cn2Q/FYCUbYphsD0DpD/VyuFvinjTHBpvVp+w9O848WJnYLT4aS3DaY
PrEOUomh8GqiVUjw45Gi+azwek3f5Qo5+53aMDCLeoh2r0pFT1Yuzj5bFKhwN/zN
wSgWf+rWTl5m1qN6vBv749AsEu2zK/sHR5GySirXnI9OvSuMrbc6/lre4HD00d7j
0vc2kH+wDCLNXzUoaCcZJ1NctUaxbVUyKh+N+ljCPNljpv/aMWwyXxTRdFpECJSR
CTfbQIkFCaPqLaEq8libbeOvdeZ/5ad5vGA16vm2ptfTqPBaAyGOZzMmuMr80zzv
B1eHjXEofMC+TCgz1Oy471BSYvWXcZyMK3XeLxGznVSTvm47sMHQdWnAbl+bjN/A
OTE+KtZ98ynjrP1K9dapwH0AzN82IArOMG2IDckBsaHQEqF0DWjxTLAES0PFMKlw
FAGU6rj4MESHUKuCc4vHL+8uI34BhDyAq/QZO7mTfoDfXGgQw2yH1gTboPSKNCYl
VqhM+AFnovQp5sqQr6I6uL3zSXW/Vgo9q61woVQ20cFzVPPwfNrJgyTYv3vjRJgt
60DExy0ci+4qdLzuzH5DJRORFLiTi8omi3woLms7YEzjpottxMuntb61tTx2LH+6
GD4abKaaG/WjMHkOD3zVt+dZnCT4VKGGG4u+Az6ROb8BnubP0aqDQ5RDDDHkdIDM
F+wUHkXQoIoTAJPbwRaeCm00W8RUM/2lICi5jW+xwl0H/DWgKTCeDKf3N1DhMcnq
rpFQY6zHkVugKOgHWajmDdJdki2ERXrdlYfnXW5BpuqM1gmKdidg1U+HQP0kBFGt
uCKUgWo4Zsp7+/vobnQv6TUO0AFFD/oQppEPuJ73gV2u2fes/ajsOWag1SipD/GI
tjyoS6vLjo+E01+HSWAjGBYn4u+u6Kl5XkqsWTjrfyYXZ5S+Akzseh3jjUSIwGK/
KAdcmivgcT3GPokUUiuq5jsxwT7TdhcDOVejL8kVjDOpgzi5I2BopEkeZkazmAM+
eXX4DAIlSa/O9cdKc2I+eIoVvOn4piwSh+KdGdIfH3LYEByaGtdRUUXh5WS8cAkK
FDkeYkbcl4u9oqLDzvE0ELxCtLetdCeO7bnwiSqjqTf5J7Vt9TAo3hhx5OH3trxm
AuDJJRpqs6D58JkiODM+/dLpCN/n9pgwF+nPyU8P10wDhn1xcGFwWuwXLh5IjRwm
8Xl1aLh2sUivHZlvkW+30vwDYp7Q+lI8yobbGEx8HhFPrp41UrEBI+y/tb9dkQ2h
iqPCC09Ryxg4FQryicKcMVS9IbW9o35PB2J20z1SceBO5JKqJ3CRszybJqh1VM33
50vui7CsnfsKMch/u1aptykhCOn6v2Keyd4U5oM/rWjlWkB+yiuxMSYd4LyuPUkp
URzOSjzfscugHQUccn8WvBsiajq0q1va+OFoCj4eWBMy2yrbt/QVBHvKQwD0KHTQ
5XRRDbkxFc1E3eDw4fYhRoikuXp74Ke67JXwl8ywpM0zlVW0rz+41IvxtFa0h07R
u2V/jp/UbrcaErfoWA/btto0eN12riA8/z/3U4SDQ9slm81EpNCeenLye9U7u0tT
LaxaVm9skxtcTUDpFXpQdrnWXPbRPL8V/hOp4Gwb4eoTv005X2iFOf6AyK7L/MAE
4uK6qm/PZSQCWS56Xpi0VF0AEsQXTuiQMmHMoxTt7bU9943Ztan5l9IhzRX9PHxd
vlo/nIerxZBaSNPQBZrR/obE5qM9yd6SOmwhUD3TOK8AGFETXSVHJTCcTV7QopB3
GUiXoQ85boOg3xKcoJxULBwBzXrQsoUaLTU2UaxzLLNPaG9TH0EXyQQBzGX5vojo
PCPG1ytM7d9muVX+b64QmJ8INSJY+96bHeISHPh05AY+GzKgdtMUV3b5CdMXVa44
FvRMsdwiBx8eme6HKFAUo+ewPy7Fri9oyPF1T1u3wzCTFrWt66KJ5fYpT3tJ2ueF
B32LkEpjDaKUn20SHmOwCQRtw2x/OQcdWG+Slr8aX3d1Ct/dK4ekFS2K9ApZkxwv
Tedf7mmVXUO8aXmmvv2yPzdyDep4d2I6FVtuRfQjh8j3dl7SkqY2CB5zK1G84Wdo
bY2eF+3LDMnpwibHb/Alko2cRQzoCGl1c+CcR/mV8L96YZeRX3CUlLDDavoSMNUa
+eom9xQ0RxCYHTmvsOhGlgqm4vlaOhTltBj5yWCwTjNSaQH3eDekzeqTRf2qNsNx
CrTHskIXH5b26BOIxeh+jzTk1m0ZbXQ3eE+YGmLz40Sds4hIG5LAvgkjtXu16/s8
vT1lgwdY4VmRlNcs41yHmoUa/bVjHW06FhcybVWmKhbxeKSIyuA40y0n6mNqFQwb
fr+tsgigRMvU+TH1t2O80PHAIb8AyDMGtMPAJ0InL6t2iK5/ekA5DFh60QTTbmNP
J0Wjw2XAedICoOdXVePASWkGDc8vHeQookVWeUFZ+Hf+eJoG5hczUFMFoLGtNEWw
sPZg1ZpYskDSjgDfBD9I29tsz2ZvQoPHKrKbKLGJF1NhTBk9RIaiVXHVqrJNdwCg
a+eU/edKcq+HHBkd+XTgdSdKw88oVBVyP+qVSZV89n5gBF4AMQsvDeZyaDsQrAYz
5V4B1VcOMoL4KUS7V2a0f5uabpdBDSTNkDt0HzMZ7JsiDQX/30Hg5+jw/UUoMNYp
34gDkT+4DKJaiYNJcT79dBx1TDm5gfgdS5Q0NVF9YFmW3DdYt7RRby3lsHwfafyW
7YKAgjKyysOXOp8bmpnLUqe/quDWLSdbml2bQiT/72/5WvtqaCpJZ/ftyavM8rKZ
tplDwBkkwcX3mmJGkL+X3rKhzwpg4JWIFofIqS4cSMgOWY/PTDY1XbS/hkv67tO1
gEign65EqWpcuX5w2jZAC5TmeChakoPVF7vaIja5VLKCh4IaLd+yRKe1L2RuNq+x
n6hiLBVlXZUDxGTDgqIA1Xc+/xGJ02E784JxJ/EqMgwCD1hnuaUsKhAWYl+jfSdA
MVBRnwVcEHhp4PlT8oZ/dfRa5ZAUar8fTyGGV04tgNqFiAxoDE6Mr574ysWRA2Gv
h4rujup/7ApyuAx5R1UYEk/B9FR3LU9oPY4A3IE/bcuBK+aNTUYuz5DBjOOD7+b6
yjLkisTN2Ibj1ZEah9Aq20pwB1wZCH9SF2B1bRJoULuM0nYE6YWweH/nvtgzAJny
v3nKjC8y0jjxp1Q0dnbTEH7JBC6H4Ws/O1AsQpTqCje+0mrb0TuODmtvWW7bmHNk
rpGiLStB02JceenRTdAK01IOgiaYop+Tm6fT7RH0MaoooALkWqD9mDv6HBfUvpEm
egfeo2UViv9PmAuC4Q/wsByJlQYERMUvfhBHRup502u+q/K5krft/MQFxxuDSwOb
lKTKQWyjP2+aKoMI9cls5FvyjijctHlt3qngvv6Yyceh8CC0ITx60I9Gmwl0dQil
S6pSVKbHeO3sgxY4YSDJhK7TwncSMxAwjNTWA6ZSpYW53F+sIJBnxatLtF4oCsr8
R8Fde4HSHI43V7wb3JCuUbcj5odAFjq374iS9fnbDdidfNqC4ZfFtyhxSuBdO6+m
ipacVlb9N4elrXn1qKHW12sJOlEdlhFyBinB0puxBF6Cuy3V36CpINbtlusT4MjQ
DZUg+nwkJKunmcTIcA0ysVQU3LwaICoeBFosXsMtx/iGYVwYAAZopl7/ERU4Wztl
SIbM8cNyTN3W3zfRwBnEEGsD+3hNUzlSef0m750ySmYu2GSEwMzOfdrMG/uA0NVu
TuG+ostF9RgUUn6GGs6yLmD3zT9L0NTJubDSjD/vLurT7sZciH4MkrAlx/Pn290B
N6IJJ+NKKXxBhrByd1gOXq9ncVpV4WuB8u2n30BsDSOsUs2e+KPkQlVVhcCE2+fB
iJTzNXFcRiW8UUEuzijZPYiniU9gaNFeB6MY09CrP0b1yeO2MD4ckonel6ctpwuK
KrEHdduoUNkHGbwkNy7EhagtIQwNSPefxF23Ez78z7t3Z5beicJv7BtHFDU+zJkR
CAIxDLqDs8CkVnBVn1VVv6hxBmjHDpkFLj1/S+rZnLYmbLtA5fC7bXY26oTdy+8y
oNJTOfp9GHWwN5lsKXbWLWa3BZiKHc3LmKaNLf4bIme1MCR2nZLxmpYLB1kPMJSG
EwHE/slFusm4WRgici2S1a6OZz2vLABHgRtHbn90OFlwfadzbSDVLswL9vxS6imu
g8nYTv776IaKdJD5uneX+JjGYB8p6FEA14F9OXm37sef3sm2m1i4EMatFpXoXsek
hDhqy9dD0aSm4WPDJl3Hfl1ciOsbwkOpvJVayRJcqviSfRTcKq9Es9/v9wgHQ6XF
MeOKXOaI5F/Au/bpIp99VOgMxVXnQmOPMpArdxRT6DAKdPxy2KmQleU1jUbdmypL
tEcg2LCJO9Gfm9UTgTMIXBWWmjVDjAYaquTAP2BmNwtVVlAk3NETDERyM51T+rLd
A/kbkyLBzk+x5Dj740sYzV8iWNiV73Nts13gIrisuX98Kd1mxrMjsJH4q1i1r6Cg
ynEu8MOoEtyMZkqzDdL2neGFAQ+t2Z0X1982xj0uOtPNt8fLQroB3xiguoe2gzCY
bhVxSe0MARnojUa/pgGkL1ox4ysfjq9DUVTb/znxAivzLJcAfC7wgdItnS/OC2MR
h1auN2pwWLnAfgDToalpx3PQnY3dP2/Om+QwFn74ntRGKenjO86PhByWR2ytmUth
8J/mQNZplGJO/k5g4wbEu5LwAXniW1eUh4rWKHFIEBNu6cYE6BfgtYhZY+yebVG1
c19QxbU3/wR9GefIflIKjVSaj1E+5XUnAVCTzTMiI1u3nKAw3L7o4KgXJ5/hlvn9
gOBKbEMgRxwiqxZbl+0AhCQrIi9KPihDv+yZ9K3nj43hGX7B+ujyy+KJ5ZH+mRmB
4qCrEOeZPFCYhP6d7w2Sn2sZdI+kHlxVkrWx94b/rJVIodZkfGxr4SeZzjtwf+mn
sl+XG19UtAWyA/ijVan30Y8QxiR4yqdSHRkqB2tlw9GMBzj0YA0B/yg6oLri8PoR
5ZLzSs3KmG5KjfdZU6sLDw76dFIGWO86D/LlYak8rcmEwf5hXdq2uEgZPiJBijDx
OxiFlK6eoGKaa28a2ygTQZB8jXfF4KlsrG0jhMKmr5DFtAuXyCH6S+Tiuxo6rw2d
mMoQiMSW4gt/1BprEug2oRWHnagkzK1vy/9EkFQuwUlHuIUPRjasolmh/pS1WxJt
cIIyERxVytvU0G2uYWKfvoohj/gcvMk7/xAI9LyvFT32j6x2lvvR9IfsJJkasA/o
gZOYhFNqsKONFuqG0oSAUfxcPHyx/cTUWOR+GWO4tU6UwRHYDDUj8+awQXCIZRcU
5PpPqgVc/m4FK2weniPRLb7Nr4vFpn2TYcOYPOvkZs2ozersHAsOSrwsvb3ZGptC
31udXZEhw3/o+X+RHyscFUUD1hGMIKPy58rYlbDhLNJMrhh/O9A1cB4ZZdl/Wnt2
/DfQcYQ4f63HgGmyTUbZE9V6JwEzMf8rXxAEblcibRR+3VeEdtNtEkFUUtgQ5FEW
2HD6DdDcYZVZCtZ4Oyqwq55I+FNb257WOQrvHYzvmTAHl+3KxStlhE3aiANDgBDo
cgZIg2gBDNu9JwJ0Peuupe8ukT1lzi0diYaSQiWYxH8PY2px68VtxaJYzxjn4rC1
hy8KDw1Zaa2z2fVn4NRLtRPV7CqLmsWsrTgMzaaVC9Ddzy1aZa7OuK4M7RWFEJrb
4sO5DIOhKRPQ+hC9+vg+s8l7ulBZLihho0bA5Uuo90X0uH2gxc2SE6LTSnSwxKXY
M6ySLPF6bGY+PaLGsC0yp9shPwpR0orWfaaaB08O6HSEbW6o1eTeK5HuxlmjOkBJ
Qvim12NHiPvUh9az96ZY+NFR4x6qG/HceXPvxukTfO54J1gEvzbvgRymk8zOVSlM
ZQl51IdgD6SdUrrn1ihUeYPjX2smhDAnGXOxwNDRU0p2xUIPoOnbMv/tQOD1yeQq
n7W7478KIFH+kygFf5p2e2+iHfWkJ+M+MWWOppUkAzmC1OUzUY0YGxHC5HOJXUle
E6lKqUPYjeAGOwS6+WDKw1Yx4pV6haS4ZepBQ0H3W9AARy7ei7DIdW5coNovEo08
gByYExjoZvgb0ZrHwSTPoXa6aaaHoEZzfMVhMyi4J7+03TQyl4kc1PsuGH4aLvub
51tM9uxxMcMfnoxvQTZSUBroWJpFgzvDG0pr9Nj6xbrAFLeAv33hCep0hl4fs5XW
udBj1BML4ckG5M+39IIqW/e7VjK18V92earLAYKHOZN39zqprL7AZ1ZBYyopAdPy
xDjMC396SFmYV/fKL3PW/TUlGuxOQokEOwaBmHD/tS8AqfNLNbzjFWC77cjysAAu
TvDYiZ1gZIGN9/+HKovzLE8Lf8l2lylBqAZP/wsZSbrq32+jNoJ5rADJP/GVr58j
nKDS895vrYeeJZiH/OfJtMllRmzrLFp1itvkarfuc5hnBMAE4zoIQXQDQB5YJmEf
gcSmcD0MMBBB+RR1Zi6x09PDzp1fDh9NcmToptXBa+IEP5ZGvuddIuZ8tyfa3SqU
DL4z1CTOxCUIxrfF2PPOHAwfoTNjGMhmF1oUKwQc0Z3rZc0zOfhkld501a6NkqnE
9HzIxAoHW1af7muvoIJ3iq1AGSNzNs6TWWwHNnGwTDwurNLLqZ2PfX//WkgCEPrC
hdHEhAMUPIcqNwKf2gAT1564f/qIyYvzo4E0y2wY0NlgpkLCPf4ZR+DqT2LC8C7f
8iKBeAeciUyh2Xe90A1HQuibqmyKifKts4DILYFZ15jUhRUXeUj+VrRD1W0tqS5/
5e6dvaPfara4jG5ivM33E9pHxr5t6WYieDJAdS5DrelKQO0K343LG3uYkilQdG/v
J7THZH8p6CB70nTY/cCwa9e0GH61u/B616+2VozutQFKXW/oUX3WzeCRuoEPcgzU
AN0f3fCG1B+f0ihyxzcW1t70u+g0UcUfICHHsSr2zFaWJ+aM4hy51gae2Ma2JCnW
TYSOLX7L3qjYh+avYJvbOB0D0PINMPCXoT2rxaO7s0uJwVjMTriw5yj3uzSDAUK2
Jj3Hu5zscu0FsQSPmCb3AzDZdSG91UXO+sGESv3HYTgEAElRsT2t88fUkrHF6DqD
W1RptEVwC5lWGMz+7CwFfVrX+VKCN6BsQ4z9IAabijev59AKyNBhbyNGfZ8DL1uu
OX2FXCtBVkrMNsIXxNVv+VJWucCYysN57MxR2AjjnBhyxu4BQdvn4LK13dcXSICY
f8pP0H5jKhvmaqwiCBJ+mSTOsK4s6TQqgkwJ8x3A1OLnjaBLxC1w6ciMYRn+42PE
rvUxeV7SEBH1l6Cw8C4TZmLsHg3m5hrx1BTscuEkJxBugq8bBsIHH/wD2fLPfM01
MA4xEIiJGrZRFI/0uquzYqSEQk4msWXMY6VYd/BjyxENYAo9N2yUMq5vLw9qrQ7B
aCJbkzlf33juvOb2SyOXTCj3qdmwbBWbuS0YzsfVvcgKMEFzlcDvEadPLWF3G5dF
yPWbLWfs/8RTJPS4uddbPUZpUYvp45HW+I8h7IwxsDcxE4kJ+lCJTsJQere0mcAE
RHekY4xEL4yDKoZ8cEiHnHKct/I/YQ7xoR1xKC0zgrxXzW8JIbP2Hs0P3bNF9TcL
HZBLuYap3ahz/00QiFsnQYOOzXg29fkVAw9Ad6DLfAorumlJjgW1BJ0lnE3ExpuQ
X96rXTkBW4/9oVWhO5mhmwgPWCoribNo20KKizQauP8KO64Jq/IV2vu8q1z+GhTW
85LeOHAkjGdOYZkGXTFF/RRbyipdQvXt7ipBHG/KbGYRby/KY7zuPZ0DS6tH9Ztb
NKxXq1c1I1UATxlWlKuYmr9sSfSLZVZ4vYDAhlk+u1KqhldEfljeeftf8w+Lj0nH
8E/aZt7nLf1MUkcw8SKBj03RlyMFgkq/YreUMv6s3ygRuVOyo8KWPQKjcTW5jHNu
NIn8NN9NCrSM0sb8Ict+NwWJtO0kTe431Gy+obiLYvvYlV7ldYGvoxL0VD7EOKr6
3/lYSZ56CWK5C/q5kpsmTSabadjph+Mzd27C9zx0drdNFtHle/YaxDOirzj8KWHW
RNJCVZ0aiLvKA8e7H8p1t56GFHmn38wW7XZ+tWX1b8YORSCMfH2yXjWf43Bj3M3F
MJfXzyzd7ghEFd8MNdTUVIW2y8l4xr5qIWk1od108xcBzMH8PWTazuYKyw7B1KIn
2cgnnvmepw53MKy3iazdTnKCOxyQ/bvdeanGdJLwaO4xyqkHXtmT6Sb4mGhFaicb
tU0xrsRl1QHpuTl1IP47BshJo7GeJ2iw/JegePwMO58oGqfWauplaBJDSE2kTozd
qQNWCmpyhdsvqf1Qh0FGnYxO2Qex5jCv5KGMzdhlXPC/Z465DGMyzz4JGXlcBJBC
f/mCkhx26QCCpHqHPoHWzKNXu8yP1JqZ98BSODcEJi+cpZKl01/DMXF7d0j0NSlI
b2Mg/SYuN4VWaR90VcVwbnNUUeH5/dXio9QHjp7NWsC0TK37KXpE4rWlo6ZYaKtQ
Eh85h/pDSpxBEBQ1GEGvzXbW5O2SmfEPPi/Kjvx/1ck213kRf6czZf5N4U1l5wuu
tvsxhNiY4svwHXqFZefKWPPPvEinWeD2Qg/kVH1FAql1SEkFGh328m1WV4FLT534
bRaapBjbrAWm2cHFDz8L4xn0RUezBlFY6d9a93nkfAXApGjplu54UwozGiOqfQDn
ECawQVcXBrJWvAU63trXUgSX4KIdsrgkuDlPn9SqfmHxFgjmOYYGnAtfVYCGVft+
DpW66Q0dnc35EtSUKbG8TsrhV5vZTV/TK0ZbLxMkRzl1+xI0VSRn0dXhoN3WBOwB
J2Powo1h5k/6LgZFyJAvrzcsKDjBJQJ8I2H2ebOtz87tmaXqLMwz5n7w8yp9U3cS
t6TAf4fwQ/OsodLGZcsyFZ7lg78Ey0+al8WofvTRsJOukSuXJ4d+8smY7aN7xnzs
jMpOtoe4fLOjODksKhgy/BUL90sUNIu4I4F/1RdthuE9gg9lqAmcuinCgcOeHUqG
WATrsyCxjrGabmgr/50rzYx/JtUYPnI2nWvLrJasv2hLyyL4Xjw8T9rHZDDOZbZ0
oCDwD50uJitdxNUdpLFx6L7Ctz7lji5jo5cS9oKCz9hpzet6UI2Z+T2yDxsc4/cV
baSwrXCT3yQ9PXsiEJ3/9Cul2geshNnEeY77H3iIlKL7da1M1SnqDFjvyQmFQbm9
2IWTVBgaoCz/L0o53dsVgtmsn4pXFd+fHyXluXMUAahygbYa5vHRSyVTk+m68Rng
zrIrYCZKmoL619ZhJAwDGEYqQPN0fkckyIYn+fO9+Tu7Ud+PCKzUCC/sG95nORXt
oI2loUb6F/QucYdn6PlEE291hx2X1EuIx0UiUu3c3VZjOyuXJHrGPIiNe7Uzoey9
LDAZ0b59/7nfmFFvIlh2AcZL/YeLnTMR3mNGn4GC4crCc+mR+rxb6mjhTzN6TapC
TVvaBatmjXVPrWan6ilkYSnXvDVwiLW7yXrB1656lyqxmmoq9AaIVf8GPe6Iouag
SgbRpXn0E84IiRG6zMM9tPHrdAsNyJ5NgIRHRnO6Ob0+pn26MyXABEsZtmb0GVYB
/JXfiOUxL3QTBpM0wqrqvLdPXMGZSkb+kLUrWv2AwHhaumfUI2p687KrxXTLx8oK
2XWGMG2ujKmGQ85ylMJTFSgOIkZu4UBrK0yySzN4S3WNOUrx0qxfl+zf2Xc15BHM
kc4HsNU8INaPnD/4kR4pu3BDwTkmSV26alR+hejl2/0nVePRAAfKKj2JeR7nji7q
hOWsB0UsBMQsDJ9krbSax9L12ITGPeEI4vAR7LFU27VqhFnG73TG4l5Ac562P8i5
dybeXcmbUVgetHcYbcgMal5aTUFI5LukfhmCk4fMRhlenHfHnQJ0ekfCDg8Pdzya
JBlSmZhszpwl4gQXtStmV3E3klSZoCBK+V+uFQBEoqad873w0QhfHLhHq22o4+1Q
4bSrADPwLQP4+FtQ8A+U4ipxTSdS8XRPcoa4Qh1Syjhf7qtFTYKmTHjDNlek5t40
tIpBqImE294wIzznP1i41jHXgQvOAnZWT73+tW9QxEgXwqDO1o3F/lpejWnHJH6R
2revBFqJPOAdtQQ6E01Z4YcJO4Aou5QkeH22XTblp+Sdgrc1v3h9TFBwDIOUXp9j
ZwiU9IJuAtPverR7lVpKQtvt03xB3h28o6IZID74Vj+rfzBAngUWJqtW+yzzaONy
JY7mgHOtBYXsJJgGFHlaeRtFwfKtsLfpSwoPsn19ngiCBavLuASnJc85c2ag8OvS
wYsyu8My6CnWRtkirgPgey4rG0IhEzc1Eq1kWqeZIEgsL4F52PEK8QC+iWsuGrko
yl2nR1nrLqnqQmJaW9g3wY1M+C3PGl0PxOXeEXPKjGMWTBl66we5I4Ugxzarbzeu
DoJInx7SL+9ASSdxp/jQohjR2TgUfz30mi/Xz9AMetOS3+tol0t1PX4Qh9aFr5cy
uMLEFWu/5aTDX2IYeGCzlE5dlDKeQKuX2v4bnWGFnbG5pBuZ1wY+lkt6gEC2gahi
f1+0kuYV2QIzfobrsB1N8UKEx8iMFguJdh1T2tkcVTo48TDZTmDJz45rYkT9dCAm
nX3hTUA8+mdn05NMTtFWqxuEn4OPZkkhRGtz7yxtRTn1qDolR4aZTdPEFKwyJeNM
X82dK8LKi5eMaTnBc+BPXbswtoSjtzDQ5D6nKXEHSezBzRsSGn19jaHcTeKVS/QC
ty0VBoYICgDrtp9An04mmzp/YwXvS3oZ92WnjDY5pnNS6c65awEiM5wbzrAbpr6h
cgoMc3vNpPbnlMhXrn4X4e/SKI8RKyJf8NHgfhUM5Y2iBXCa3ZzILQyYawApmc+q
29Zx/8CWd3OQdiE9t8UUC8rhD1Fo0wq7k+CWZkjcwRGolfjBt7wRY6ip52ahACBZ
u/yph3U/v3HXAixZvw41DmVrHEaJu7wuxl76GfaxJncxzKFLJNUDPZEADxbLJGqk
5UHj5KVie0a1cwaEks7BWozN/RXs7Qlj+SaEyZsj3AekPtiV4jHINE8URko+rlwy
eKS434gY+Hd55ryeeMOjcm2d14BcEnnbZb7Ymjls5F9Pq8JftORjwAUzIT/hQQQp
dcCpq0E7vxuSLIs9DhqNGW4fC569zDIWlmUHgNxLwrIIDD3CR7TO+acE+tKEw8wM
0UqegedNSyi9PbmRvMtyO5M/iaha3fNaVMnfeXzCrwdTYhWzMFd5N9KTQTpQW1Q8
Eh3WPg5r5LAVsynRnC1OueafUodH1wGePuqTgaVMxpCJCxhZaGAeiZLTD19nVwi9
7lJcvgvcBUKdKERy8h3WuB3+MsQAtAuclIcysLaL8HtRjiYrVyPjbpd2C6Mahhf0
jUDXneTfOn5lV0r3anpx8jNJGR5OIoAT8rKS+CRYBAnr8FaC0lo8TG9XwE5ZIfLx
Uit4whA2mg5xYqE/qNeOQCvXa/A5eIAQsG8idSMV/5B5z4//pFpgbO+V1/YvxpGS
O75uEm1DDu/invq6YYgSHsqBkIv6vpT9mJv7kDukas29zyCck4P1uDz1D9Sg0QbR
J3ja5HB4L4y8S1uOrBaxgL7uTCDiI0cYGr50zYV5VzlftlfpGaC4MXepe1kD1qCk
umIJ+97K2JojM5oeO4hZr7o59Cp8PL6sjpVcRje2d4qEf8f1x836ksGvMD6LLLF3
yvx3tdimajIQPEs44EBFF2mF2s9jUjWx6Gt3bjE/h9m/kJLhvvWlPmOJz3RyZmCH
zsK99KeFKPb1cZWYHXSVO0jMUdkf9s8s/kl1uK1oxrU4XOM6mZLsFbFORi8onJXW
7PmGwNEdt/g/LyJqJOu0yiXJxD7yu8FPB7ZRgfYNYBqc1eO3udhuYqeU0iMLgcxv
s1/R6d1e3pCrAwvJjC4pyxyZmVnaFhNaaskg0N8YqHsQhGgDZmCJYRPP/I2vcilf
/7cszzPrJyas+2r8Ufkkzm5ug5kKEj7/zSe7z/2S7a+hFIN+rnGxmrbcTU4sTMFA
hBZklfLUSaqjG+TsOlLSutM+Z/fJSMr2SuelT3znObNl/YhN1/fvp4icLsuU3Ry/
q/eseLmVnSO3z8s2dRPPFptOG+p8veMuTacXiLQFh9MPcwRvoX53mqvJ0d/WBVXz
9v/yHHBMSpuQyFTRkKa5psFD5TURng1ZrXNz0HmtkANxeEdwhv+jnjL/gd/+OgGs
twcgjH+jFQfCMFQMbtDFwm6H34A/qIMEiEGo1qOYyQNYA9xYPRQ64imK/3Sk6DCm
XPpczhOLJCiIG0ONDWiv6NZ3/KL6qqkxA602hSX+oWMvm2Snns/5l3HYaqlp07XU
I0kqDkafEo/000NsBiDPvTSJWs8sReIN3PcJEfxA/WGuZ9TMzzJ7zBaLLSHv2Dwr
3oGY9zB85wUz5/uJYzJJCCiaS227AAfwZxCjyDmvsxt/LIq18n2QMYIBP/z64Efj
SaHbaCQDLYzqMy6Qkt4iTVB6VgH0qBTvGocEQHyUI3TBwa4W7LUAoZ1wRUfns5E/
TRUfoahbk/0/vS7CvCRlqJGsJk3kgisWL6/6UIN7/TLVwYMXQ5VRsvuol055U1cm
jTqbe4Us88lYWXwLmGEfRggkjEkUHc7k5If5gpw5WGeDRi7aBP25xEqFvh/Tcs77
TzwssJg1tJ8OTMld4KBWjqM4cYoCpWsvzzUDasAU/hutGlrE7sWNrPViyrztd6P2
7Mq3Fn1fEJyvmeIXFJy5NfBAr8kfqvSlvNoxwZr717F0pOTDvsbpZKAOBjL3zEiS
OyVXBu/s2dT5bNwTeOCFvCQwNPoDCTMTJRCR6IV9GrtihOvxnaWsPyKOQr3yBEjG
Hm7jgSR+/2/HsQQmEyQyZKlNx2TXPe9f0jO4mmiCihI6hVhjKJsU6ciZ6GLHntZH
a+cx/hoqE+rlYmDAK8teK7qXYrJTSiWImqRlK/Lkts9Q21qbC7Tw8XquC8mVMnAs
SKl0uIYlWw0Rmu+UunO43VukElnJi94UG4kCML9/vSKOU3aOSPimRke+nSaKqAnO
ZYesjKyREawPdiHWfiKcC9qu/OlxTUk2lgQSjvI0Js/JTzv/mi/mI+hlqFqMCFNr
cCXx2TbnGSNqbsucyFwNmOXNPPRWOml3P78wvYw+UpBu15Uuh2y2Qt6kMkGGcinL
Nd16dsBDBVwWQEyDnVWHWlel4LW2crh6e+rekDv0FWalFQgAuPrevGoC3m4Vj6V/
CepT13i3nh/JOp/8bY9lyX+ZAcAgBIiPFF9E4+tFtBPLSsqzKJ7KKUU0xc5+T8a5
j73rlw3d6TXjqKUBq7BMf5Ytqv/3++RjuPp8656ey/e8M0D0sRfEK0ndR1JP+ECa
PCc2XM79Q0N/Evh+7A1zTQDhGgsdrd0ExtirxSqnmBIc7Fo9PzDKum+Gkck9qY3H
GsP5MRN380uf06511RxkTeBEcV2XIKV8qWqmJTFQ67/LuOQhEshRkOODhR4jes2x
k81WiNW+z5lZpixODP513FprywVPGiRMCqMtsAI/u4BxXPuy9Zc/oSeTF8Oh7RzL
9a9PgJYBYeMYJvk2D57s4irFcG5n0GcZBrhvvzSNLammchEbD4Y+kzaethCAA7Eq
8jfqq7dGYVs1UIly+DX/VFFZIjW9UIglA2GfErf9/DQuOnYHjX41eS63MIRuk/Cr
vUPDH7Y/+v4hDvjwGAB0pxn0TdtGtbQmO5ILzrxTJdWkU4zJ4CxJTiZ7xxlvgi28
sUVB8j4XZE6o4S9DDfmiQn+vwCBB8A1sP1vA3OTm+lCDb3yhM22rsBvPx1egEC65
ZD0TZNa5dQIwhuc0kFSPb1KxqLljGZG3rLurCpMeCFGzA/tPaEgJLUj5EIyKs+RT
h0SYzKA2dguEU/wzgCKXHYp756GgtNCDPxfrvAAEtCdnCBP/hGZvc9c6wN87vp6D
OJnWe+HuSqlec79wh8Fk5qOcNNaFLp6ciDbgidIR8uY5dyHef3TEedXoJirVAvvo
WPuMy3qengDIoXnigbDkp+82IpLOHb0O4WvDGVlzDcndiuHLHXk5/3o5Ssh72gzh
abiMjeHr2XOmzCkjNV1XlTJXpsdsz8BJTyv5hf/6PwQRz+exbJg0eETQGYm0aQJ4
hb2/2elFFtePhp4g1bfFFMqaaE95O04eGwk1XszzREqLG+H2IYnpnbO5K6H/wwf3
+8WxpO3Ih1IWdb4g8GYALQKrqzkQuBZs1K8E95kSiYoTYRsAqJDzKfDZAgZl8Nzd
8SiQlVvA8V56yLOq8U4a2Za+XCntNY5xoI6t2iWLty4YfZkN4FthL2obt114dr/E
xbV/OS6yXM2bj3GP4m39936X2siKBAg+pfw4rJ3ltb8aFKWv/F9RL6G2qGgXx9I2
tpDogwDk1DbEngMFhGScI13JJ5sozeN6xpWYMB/34zzCnW1JRRk3FBG8xSvoOxDi
FBp4Hqe3H/pBHhLUVd9WdVW3vFttZlAo59tB21bc1EQpqV7VtuZ2QuczIamjVw/q
P/LbrQZ2XMXIhddFCSi17ZIA2nUucQpOIU1KuZEZPUw9BnSLfBOWkQYvPfwI70Vh
3t630JqO5+nP2x336ocQIfhJ0AbXaudTvllcIGBVMfD2M2VAj0h5ilZr5S5gXYGr
IuZZG4YSOMd18y2Kzqk0tmQM+5DW/H80/HtkvRoQh3XMts+tH8LhwRfOtxFXs77m
j9rAJlZeNmhVIgmb73Aih+w6KRWV6nC/YY5bBVT9ir0ddHArHKK4nqVYW23AVQtO
PfFIVChgXr01ZhU2M4FZbxxTVHci6Okeh60njy/opdpMxedhK6W8jJGKh/FLV6kZ
2Ac/qsxi/RUsNmBEnWV5JRM40TB1F6azYVRBjBFssR7BU41g06AcVPZTGdAEYmfZ
6THu/tv+WZTDMhqem8Hert6wNd+8IPW2NhWJjdsBehS4J9sTjPAmeNFQS8mgCBb2
ZDmHcKWjE9bLqWNyg0rd477BNzd20TBP4kmKO+i7wlQuCBbEu8fGTby6P/lGrqeC
WOw9YbY7aNnIqFtJHKxC7xdli6n23XJ/CvoBKrw8fOueeIW/71jGEypAi7IClWVZ
jxzGT7X17EnXErmyW/a3/RUhcQsHGLrpIzDTGsXsWP2+fQnh4jhGJF2p/EpF0ZJW
9VE1ud0bpAN+9zUXuRDNRNtG8ApiSuiwSZ2vO3xPUpNogiRWS/BkZjgqvrCGB/BT
QWi3lJKOB/bCfgq4rywPR0gU6uqVjIk0m8swDAPkueV4KURaGzJ69jwhl6UFNGG6
0JEHdJE6hJzdIKIlFJOTDqrqEXCaJEV37JQbxqHNQSupof5N+lb4hDpeUsZWY8JC
mUuMVqJqwvlkMkvkaSlpREf5LjZOYnNJNJDFhvBu3P1vOa8smSWUbUkkragRdbyv
EjQsVebwB8AVaxpzmt+g341XzUDAI62G5PfdO/+TwyNgC79Ldsp+h5ARwkQJ0gLY
Mz5MnMOqpJtYkbYHU38amm6aEWLYmArWWxSOqBU+tWZ0gjOoMkYjVFJnUl+KWXtO
GWp6Mg2rYMtSx70yM54BqXI7bRkI8lPxd6wsSRSJkFa9mxgdH3VD12kl/xJjTJx5
v7kgl1XIwMy3csJKrBxzYmWt8f6kdhh+9IPCHZxtd7md5aaxNsU5HphtKpqgNHV0
e/qQ/1Qp0EpoMq95f4LjSr45WnLrfIu3+VwKFujN7pEmE7HhFzFEKyG4VIm5f2ma
8jPGUHc/wf++Ms27DsFg9CKKZCpfmnBjrT45TFKvgv75Rb2jScTtYPuAuc4AxE8c
6VPg5ZQ4EDmZJfi7/9RWqVHWuY6rF1Ce+civwJNoWpak+899JMmqio29VNnWPfDH
g1yDX+C97blLbysvSOtsHfR1SkrYZgpXwTTNoCkvqtZNUf8xfP2x/58xu2n2QxMc
aJNUnARnCy18Jb/rIxw8oEMEXTn+o+F1L2Ji+AaVWjlhZpcsNmUSyWu/qgH+cHvG
l5AkBosbVNcuDTQOZe+W3assxVIkUH6DmQYk4SKSDEEkkJa66K9MySY6AVLxFROr
dhCUTVkdWy8XzRJYi7uQ8CZjITssYyWrq61MVjBJIpmXpu1gbTOTo+XKkiheUekb
SaTjzC1s4igqzNYCKEknigZcMp0+yXoiXGMe/vB4vsriX0amkDr3NPydBxOKcGUo
fQU4PanYkDqWfM7fiIfHZcy99slIuZ+xXCIsr1wczqxMblpZJy6OQncpYu7CrjLp
OXEFc9uStY077c9S8vgNnCvPmnKmRYzU/ihxq7C8IF/5VCeAhcvIYgBXQ8+LiFlh
tno7QOo/ImcugxZK8d+qDK8RIG51zVKOL2MFmPhLW/KBl8PIpGPlGFOiwkAKPeLA
bqjtFUep1j2gEk2GZdsqx9jKfJ1I9xYur21+WF1s0ZYwbc1j8Vg2s6h2/YTmHezY
hQJ9wUAEn1AzHUOQpm3T2TliW8FjpuQU1FnboLRukZTzyEpP2dw9uvgrZdo2iJ5g
I8mZsaaP8cK+++L8PRnQ7XuPQvDPi+DCHyJHl3Mlvzb9F8PCXfN7vQQ9ON3lQigC
mnNIfXTCn+q5ynCyEQz7zjmBAdPD/fDZe/kk2bBopO4CqF0Kx4l0PD44DB5OE00n
LkTLakFxhThcg8ehU+O8EEvNcTILtcs3yAIYF6Oday9s2oO6I8mZRUxIQ7ebVtM8
kmVqTrK9xm+fvz/R6j2ZJX4wVEIElSbSeCtGXq7x9ZjAyg8omX6LWYyc56fVrQA3
gGgCn4XAv6X/ygmAB6WB9aWE8uwQN1avN+Mq18fz+EzDADqZLddRy/uIn+Ne+5vP
wt+sX4b51mymK8KYjpjGE1UgVUPJmmGz+TK6gRUmHNE5eaNeZer0HvnGcU9avRAK
Pv3IQagcKh+Svnnvoz/x6BiN/oLXeTXCmjE7KptQ3X/TgcwBd3YEA+gCNkAlQRfW
fs/o811PAqEF+oJXTRe+RKoehqDGpUmu30BDE7GBTlkTlXqiGgcCzMu/lUX4tDuE
q3tSaj2WqvEC0L4sLytGXriXBc4kv5wssTmxShZDUvxvBgi9h3ZHufrIL3L8LGUw
9xBpUT22Yf0B9mrZSZ1d2DoFgKSwUvYT54T846oO71FDp2r4wbtSq76a1YFGHAK3
DSg698nBoqKK7NcaLvEwht5EFyYb2aFScNh4TdsO607xSnsqRbtHvUnfmULE5ASL
MTbHqu/2qoXyiMgxDknxZFzgxqcINmisJ5DfHT+mKgVE3OaFGCPOXqkXe2Gd5iA0
WMFH8NcA5TkeO0JUz9Zz8yKHe/6LH0cbWv2p1+nCHIPM8wY4ZG4LIOmMLbXzPObJ
OqQQJQs7ISjtSx46z0xpz4PcLgfzR/ELEqVzgONve28n3ZgDmvCzNNa6H8z81EE6
9sJQ9kA7lT5tlPEJB0OmyhJcCM0KH+ieNHBBi7izMhnlRvUn9L6SjJuaC7rzOOob
8eqSWDxMDB/BvXmk973f/zyHLM6ptkpHu0L9QNGQBaWvxoPWDG3vPkvc66t9TVfV
RefagCN15W77PwAhowwcqrsjR7tvarNYOqyiELZefmfb+TVaM7u2hgGCdSAzDMi7
/TtKFcp4SCte/cV9/zM5r77XrVoePhYoa7WcRvUOf/v5pxH/h//QZ9J6vUO5Ubrn
74M93J05HC1ys5WBqgVhPaaYn1xIeNyEdBuTfx3nfD9Wbq7ZfkRSRcdedF7WbBen
g7igv56pspXUBDQ/PQ2z8KqOq0zlmul9L7LArKURakUV+t7kQ7NVYKcoQlmNGPTO
H985iUQNspKclTfgUWEIEU7nn4kvVbvTkrT9xZuA6q/pqmC5mDMnH4aRTElq4nNT
VTdWNNZxBYXR+Tk2+cBI220iD6TDxMbD588yVX43wIlIo+C+v51ed6cuTXuQBUhL
kyppGUlozERDCMJDby9VH+yts3Dft36UCHULBjjivMkEG6e5S4lf4d3ucKfMetnv
B7mf/sRF1gr5++v4JwvUYiE/qH+xVos6phdtkPluKSo1V0kaS34CnsOT+CwRGi6G
dTjkpSd7r1wnJnk7BDwvaoAe1PaYO7BoRos+yyIMUfDfyNqr7twjqiFdxTAn+C3p
VCfOiIzV9CXMu6VSwsnGyjFwOiE2X/NpCfilfRT5PWSb9x82cRQepAv62B99r1Xw
nLmmP08hdh6/kYE+W4iDFbYIMZ8iakbOpN0UWPajdxomLRgjogOCKOQbZpy8GD2w
u2BhKSV9hZP6Z2DVcPYejyrtNQvhp/ScUVPToh7xQb9hcN1HrGpbPi5zNOYnbMTt
m7E5h1OFHjlWUG7OGu23i2Nl/3UBuEKcYvEndJmSijp1o7P85HFNVI146ic2DWW1
WIABJUlVkUUX08Sd0nL5lfBqKmlTLKTKbS9mgnKM2LYzcgtLBfwEaqxFOno/kC+s
AHb3NVGIp0ftQeLFP44abPeGinSAJx//hfA0V4wd5qhP/WS4CchjSSsJkLTcWje7
tw7WMR4Qx9iHGRocS32n6HNxFB9qGpduWj4YlsqGeEbSdN+Z7XhSqe4Ri0AO3WU9
0yQySlPtEC4as6OCMr7stIXtBbIhjUI3fIfHv6kZEY9XlHN9CrQ//HmR0PuIWu5w
uDkKlVwXRBe5HGWdz1qVvkt94bfdEG7ZSMbtY309hX4n5tilAuJflsgaCpjJ/x01
4qnJP7JcO444ATUVwUflwGsFbhtYFtFnV/AwF4ILO6Uwv15cqBEdIVmVydALL4mq
WBhb/NxXgul+6JzFQp/Pbrg0ISUXiHMo/QD19uLRTRxzf0FHzwouZodrDGopkktX
WaIhfWRLgTu2PrtLzE/XAwgMo1N4gYmCnmw1ls0DwLgwOISxjUTD+Q1bH6/zwNnH
tDIDZAO6uefhSsj8hM5DhQpi5xe8T8Ur9GjshSoMATlsfBHI3Z5cSWzz0taoFuAy
ExmWvWWP3tHcVH3L6Ddqh0NKyJGgu+PAk712i2EOrIh3w3cL16Mji3uUxBIl96mo
B0X+hyS10apd+Xe35g+MvDUWV1lLg7ZMGFi57wbDKwJenxx4eWaeTdIjHkDMjupg
qUYeHT1pCjSkAb33s/JXNPqzYjqOR2sLaZDxL5Q68wyehfDm9KyTnwzHNSe69Z+2
p6NjiTGOZj8g3ejIoQSI4PryF0HNChWMg/Zvd9JIM+BBUcewDA0rpaIsVxskWCxj
yOb49yWmoFE9vB02hAHRCE2GQxDB3DJOzBupnpYnrgWMaPQD742KvuuXRcm65YKO
RXRHYUPumD/4G5MUJkHTLcyJ3QbcaAxFuI2MJlrtvJ8rahSqJvnarx6sUUOXArRM
rhC6OW3f4TuH/31o5/goJR81clntwmlYT0cI3mdIeFSjIA3/aUXRrTJgrXdWI5WL
0SKF7hi7JFBcErW+gojzDbFCuyLuu5WR5uHIOJ3UOTx1fcPANsq3xIHPXILD4oJu
j2Eao0F9DK7kF9bjQADDyMcfnmoGyyYhkxGoAcXZJBImluP6cjR3QTbSZXg8dY29
EpEsArVwPBC/glW28fRR/QDouC+ckYd8r4fMkitmJjZbak87w+WRqfOmL8nqr7mi
/Qkj05nyY8ainE6awB5hbBrooJCVSnpGsucw5n43NYP5YFcoz7BAzaIwIwNgyUxu
Ux75SulQyD7FvlMejeofDPQG/0WsAGYz7HpdyviOTEC01OdW/BG8ZD+J7GhG6UUT
0Dwdyp97J64GdTrIq6jrrVs3rvwc2Md/pVY0GnTWi51kIts7GjrHsDvnrM118onr
SxUvBy/ooCFBdtu1B2MGhjNDSySlkPMotwuskXqxyCNPlgrHWrQ+gTjQ2guJYpYI
YiEFy1v3lNBcVz4VzzxmhHoWl7LCbMni/j4ldiHa12fl6fpnl7quH7Jmgq5sZEq5
oivcxqpmz8aFciVb6fKHhww5673tFaRPZiqBOOEbabtfdgqvRxAocO3mjOfrDZZd
iw4e2s7uqKRBn/B1btb7fR1wu6EsssHGpA7pK7MyXsxrprMOH9VRo/7jRww4Xozf
j7+XfQe/+uEx7fRzTCf152PVBElhOuklYM/CUm1uItbjouUOwZtBaH2IR42o2yF6
pvNXhokv9+1BAK0mIEDrP0l0mOeQVmMKuWgLx90+aI4qfos7lZ4OteSkJ9lDdLSE
eg3WsFq5gRIu4MDxUybvHXyri3vTmJXPY44BMTdxa/07DMI7FWAw/uqR5KNWP6/S
80jGX6zWczhTqEDUHK4d7aod9XoJjyYbe8P+t3VN66o+75zg2PK42OU5AFzHhXXd
h898B5KAw7/CGZhWsMPuNj87H1juSsqjSTf3G+oXJcHZzPvfIJ4yprzxTHNownQV
8yw4vAyct1bjEhWdwceSd0zx/uq5jzZHjZY9umC/21A+FU31tu35PB6QexH14Q/4
A5dTpZIYdFoM0YfA5nPtPyWhGjQN8RebmhKrlZMSgVV8z7FVQj6h9JKoA3QB2BSo
IBExhGG9pa+A+JZHYhGC3Cg1G4gF1OnG8p83ENWRlUc3lWDchkGYWU5STpdbPm8+
/aZDiIA7oKBNCGdGvT6ehbD8Ywa/IhPbsFUMqM3YpTI4ytJyAexIEctWlQUPFt/J
33HIHPP3k2Bw0HmNXuXOzu0cFKzzIrWlLF0GyFOwj00m4Br78C1IXW92z/2gGFBm
Jkgyz9Vi9a3RJnlaHTkbyLZhqsh051oAfvbgX4CpfJlB0RBff1Dy2Fc55GgQl2jA
mu3O8WAbkY6JgH40LtIDNJCnT1x9PZig7CauNWl38aALzR4abe22YkhPgLQBhqiw
iHI53r18zBgY9GKvWsChmsOitH0v19mUKDSC34JZVXHUyi4ZGHio5YG67ttbBUfL
swiMJdji+g+9mNns+I1uBcLwOB34iA1SS6WIMrjI1FKnuuwZyqL/+7Fv9nd4kFIu
EW6QADbhh+gd+HoqQKCxbgVnMlhQP8eGbJeI74IMFF+/rr8f9agbBv6wk/WFAyEe
A3Z5oCUJSEfknU8C8qg7wQCtoeH5jhN8D9LEusLAHydRiNO7ztl3wJNSf1p4hfVD
3kFzs0oOkpEhCvhV3ySLTbcH6jVc+q6x/nyNBCde2ycmy+2Jcy1a5V3UbSRXwuEd
Ptn8BJLXP8TlDyHoCYhPX/LWWcXaykJZj4nhEUUMVKsXgrCCDIE7ttR6WAzldkNn
Nmnk9RSepub2HVa8FP3bNn2/v+R2FUiDe0I6OiU1Tg6LKDI73kg72ZGqS1I9TAsY
RyUdxG8SGroZjKkLnvq4vD8vxUJ9JerqyXHs1xng0wP//Hn1IVQme7Bwo7zBJzrx
a+u/jt2s8JBxxpd0/9kYL9Fi7Na+YFEe6F+wfY2TvMxhtDVNBBZ03Q4PlMgzsjRO
wv/5INFRDYF5lKjRXfa0gB+sfyCDODIAPvcYy1zeqjbECRh1y4ZcsRakVc4hk4pO
AW0wRqdboWL2HiqL0J7zMbZwruUm+BKE7J+KqhHU2dwkdVoTGxMcdJSYCoyJgxWy
VECPavYFCNXxs0+8CqH33D2A6fng45YkE+FOoD8CKlP+NkkkWgNf7n0bh4wp4HGO
/NQm/aZtO+uZomKG9G2e51p6erm2zLsDh+kH79YkDJIeIC6dmB3SV64+a7u5UDae
25xu9x6LU+HE5imZlLeEhZTpf7Aib84g70e7Vcg3VnrwiEGETkox2OriJqIWuvJ8
BPVaEB4FUIlkFPYPkHlwioOgRj59UsqAOrD62EvQXOIwWexhKT45Qjn29RBVyZJv
U5W/CGf3y2EgZ7seEhY7bVAOmUCIK1L4b1J08ehaLkYhbz/vcU/UQKVSJzwCbi72
XZrvLBfGBJVUxBS/0JtkkZ4INM06QuuoH/JEVIMt3mq5ysWF8vKbIelHNr5tndDu
HFJJ35VFtSYI0gCPwE47+6oVIec9F8QVq2ZYs3PKw3lY2ziZhQSZDALndhfeMKTH
OSl9oIFqIgNn7tDEDWjfs/yyf952Fj863nSgx9ubyyuFrsEYVoOBRKFm2/q+iUqL
3jUukPvtpCfdkruILHridwtvCtd9EmegZ3JXWYFU95UJxI3RXrO7ITAv+s3Su10b
yGeQid4itR4/xxcRX/owAXVAHom9wKbU8DrS/ksgn8oAbcLa+u3zA2WaLRuR3Vuz
5GCe+dZKLvhu1EoqsTkJAxFrJN4Q9VQ6kQNU2TFpWJhsLCvCpfvYjOVsvIvXdArw
kkVxaVSuTCMf/z+4MurC5SqnqSq+TnSPGvnwkGcAHM93uJ49P9FKFOwWm3egwwXN
n0UzcJNb6CS0aTqAyWBb1xVo7hRj3DiTWI/QKalXTd9TX21DHKcouaDE58fc+E2/
Paik6Ap2tY4518CgueDi5qdOs8A75MHIKhK/JL+REjyPh4lBP7tHAeZjNcQwbxJS
bODv5b14IiFNLqR6iLdQnFpYOLep4rPHCUgWgZQWqIqsnzlZffUPT18kcc0Zfro/
5PNFUURItqRlfV+5G3HYGnS+0ZYkqd1cdP6E9yZvhJT207Wb6fD/ZKawcupZkiNh
EhVMVPkKs1gZ19ZwKyxSTUY+CR6PCe+T/+3NEJbmgh82yt1Vcaq6NmblEq27uZlS
cH0ouyUR63Isxy85uftmB4u5Li51AFhe5m5eOdQPj6o76lM7ACYn37eP6LcT7KxC
FdvgAqbNSuppUciJfj9UFkZ+qUKitllRVZ7ShGvIrUYCuPKSzEWu1jJvK8CqIFCT
9nLkatpb2cdRa9g9Pe7vWDA7Mp9yDhA3zK2yoC/vuTGpTuewScYS7ryT+k1d+OWg
kXNbCdz9jp9lm5QO1ycwXIoGUxpSDfCflAIZ9Ka+AX14uN8rPGs5+1E9pg4nwslC
Tu/ZWsytxpY+F0/KuVlgLDUUpeTuXW+nBq3oqwvKwDW+1Wje/O2nyJt+FLe9cyBa
5VWM0JzE9C4ZSme31MQngzJ6nwRYAyRbz6TpgL0W4A2OekfTvuNWZ0pdfDZ3IccR
zxdnIHRVAx8pXxGcweSgnGX3X+ihMH4U3C74ouVPba5xkwot2vT7z2nzJ0fxA29Q
HOfyjqY1FPC1eaNjXBp42MgVkHbH6XzkLhLBNTpz445EjwuQaGtzYMeGA9Od/J4J
2dG2okPuikhvZZqFVMywoAUeZ1Z7llfNmeatxAZuHAQMIfpWDjdw1KF0ky5OjNcr
hxBjJYwZJY7WPacnvRLlvYyyLoBXzw3G4Z5u1lJG74T1HrL/JjlzC3MSJg/4t4wN
q2J0p0Q0YDT0dtMCzJLBzBVuSr+30qQjGemZ3+CIINPghz96kLMhI/Qd3fhZNfoE
t6rtiJp4mDyel1gKPlua1oG4RxX7UphPeCJm4Ivw1ZCFLExktJDVAhFbNUod1iNq
2JAqOoLBWHOAB7VwatZKDTFiAJZygtDFG1V0BF8Vt+1/sq/MWH8DPFmjgfsSAv7s
AlrCD7B7ycO0HRj3U+rab0MekthDO+G2aEJAoHRV7+mVN8CLlGDSAM64Z85ziTra
9sxEsWXrSKOIwTkGMq4cLBJD9D1ay8XARHnKZz/JAzGip3EGdFQg1ALtBNNLBlV6
DFdjrYe75Z9NFJjnLuDTciz3Ba+SGIwxgdICpEB7gqb4Vp9a8VRreiKxw7W2VTdP
rv9d51Gjns0/lufzpqWHtfxmrJAJJ+xfm6J2Uer9l6OSWFcYI4I7070ViD7w84Ew
7gOAxZXZxEtfQabMICTmQE5Dn5duCP2ip8I8+o+5baQKVqwbOnTwPvMMAUj20XzT
zvGCV8R3cJd5lgkDzODjcIAoO5CgDfHoU9n7mb7Yb2eivsPRkLlZrTLhH7UVNqFV
PHXap2atTbNkwE//ZEsY0F+CDbJDklYMg4tQZ5X+bR94Yg2SJrvrGquko06bQqtn
Ert+uiqAtGawHstkTnBdf0nVzg6/3//2e9hFmJpwLLFwNoDRWCO86XGTZ7NX+ktG
61fZ9sttjM0FUBLFpoMvL60w0u/fD5LI0aOlB01dcevscNGcUpsnsA0XR6GWGv0T
+inT9uCwQVMa5HOddlqi1BhlO1EuKsjvExSQKeuQE07cG45MCouPZV3zfrC6mlnV
qpJF2RD4dPgv6wuU2A2KuYtPN1qextXzCB86tANzjE8noilEPphLiR1UWS2N9iD8
ja2pVZwmR4uYAlznROAFxtyrm+XgYVjSF77nbt000kMlk5RuImDSTyXHcoKadyE+
WgJ8swWcMMqVPmk99DllC+PaVuYI0rLvZEZp5iz0MhvbXn3XWGQsGsUkIpDTGCjE
Ak6FqsvZk3IkoyHcmBM++aDScSg0VO5HrZGJgog+WVznBzn5oCoQACfFA0is3dg9
kn2+f+SdaQBur98VWfoAG7KuPRtkPVVqkIV0o2w6zZYf/Q6j6UGaWRPT3DdpVBB5
xxwr9hNJ1A3W1s7EehEK8/X3twYytZajOcxMYYXn7oC+7lkld7IirxdjKUYzXzyt
ZSK5fy1LCQ7p5A9qAf6YC4u9TSMHep29ynUewx7updkxLwF9omRQjJ0qwguGzmVH
IgxrwEiVixnbM20rNuxDOLjlel7MJIv+8EUoajMsqXrQ84sH99iM2ducyz+u+/H/
wbQoz516zEsWHAhAd2SmHaaWHtKpDUlLPZ0Hz5kR/xWc7Ym0XlRvJLdrK6otdTMw
k0uhmJ01UEKxHHEO0y7w7Zse9AJZtLeD21nlMKJ9wWtCyRzsK2OJJwz6ZPbV1dqW
8Bjwe7T20z4BhYwFlQmhNhvrBXPTus7GVpND0rhaMoNYnaYNnZj0c3xL434fuBIr
+W6vrngyT6Sr5TSqHOTPREYXKdjSe6si9IzcDJBRPU7LH1+yCzLqvNyBUVnOvJlF
V/5BowyA73XkSJtDPKwfu0vkWv/9nmgfsvFSimVU5ujvtP8Z/N9YFy5f9JBga0PE
31J4vfsDFmv+7WAheFR5JoEfFwAUfHMNcy++3erbIsK4dra7PP4EgDRFlO7iR49K
nzZxGNSIpbmSnpOQqWNtI53oSTSxNwSUjrPBoRmA0/77IebvFWTLaPv5nQQH90WV
4HdMpMVPaBYvmDoAp/6IHmdxhfbRCRCkLNiSSvo61T+QSHmgu7IsL8+7Cm9vYvY3
A3jHSswC2NrvuQNoZh0TIKbs1klYmhm3zZCIFjQsmwDUC4ziIuIrvE33ga02i6ht
KOHCUXFq3K429x9nZQy9mfITgrcycQ8tJlZ2hAD4g8ajA3vR2xzRZ4JsomRnP4kN
P/jdetiqgb1R+yc5LOype3xxaQ2tTG3VGYnia36Ydg25ogTQuMZXc18SrrIbeEEp
tbhSfP+6XhIQU/RMe7054Wp1zOetp/udZJu6MiCDEWMeD7jED2kNv9I85HxmcBeG
HaHcb1YTyY1jVwuYSk580Kf8LBfWwWbUI90/bE/bBDSYT9sI4YywZwQIwmUF6BTb
bJkxy8hDinfxm+0BkOyCBUWPX2DG3MKG0phKRqgJsxUW2dkWoC9cQVaoJFnEu+oS
eIuOE23+NoylXq5xgf3Yomp3keCGMhBPceKeHhCysXtgS0kZgVU1Grd1zWPZtlTl
yp5r465/VcrvOZBtLxGC7waWClLPSk4BqgWzTyMtsSBzsjOM+W2+Wzz1GYa9LW24
fhRf/HQzAeZBRNgMUqPKyU7H4rHSFJAR03NpWDU3QEaaqbOeSJSwvTFbx5TxP/4F
ykVaPz1XFfoWVyy7h747zuaWhhGklLSYyn7xs9nKv1O9jsuInmA28UsBCrkstccp
C/xke3Cz9SzT9+Sgcr8+Uf14Ivk2ffze1cHYbRxpKxO8gVL73EUejwwOHE8hUj5m
wgjef2z59zR1JY/Sff2xIJDP7fmEnR2ysZOQsiUTW3lr0C6VUOmxWWFrUxVU1VdU
k381JTCUvSPMleBlYscRqw+ZJKuUt0z6/kzAmy6xvhv0lWqjt7Jllc7btQfKFeGW
qaZlKuBfrDKXwgFI3Wut8r8zJ4QazZeqwB8otaEEa2zrz64Rg8/oHXr87ixmuDKa
uCJGKhBntMTtZ3WIalBawsC63tda1fMg6gnlLqWe0NF5m8kZ1LGrbpfYwgrUbR/I
PLLmVH7yVL7GIdNN2hG3+6E8idwLZedkOTHIGNyMQ0Pa1W6URUIpYOwbS8INqPRQ
xVnlXEr330L99txbj2jacLZfg0yx8bPNCOPZ1ctZNkhNvTTt/Xhbp+WSx2Bt6GMr
iONI7Aw4REeAuX6XDrVSSDDnyc5GVnmPXejsCRNHJzMBQWccmjXml4/t1KZ//mW+
7KRuA2dTs9iJfeChLG1eki2qOJrLbjH9HDU42/AUTylqnrnYhGHvagRLviVweP3Q
hOB4jRTV5KpHwBeitHxqQ6O6Vpo7fqNXOZFWRwzUZu1t5V3i2WxxfY0EoB9gbKkA
3U9jHmf2fe6bSRsnTLtyVXRV6tMGT7K9EFxLjn+5pT87iyGY5yG41ImTG6GHvKVV
Gn5s4PQImHLrw4UBn1dvIVlUn6O067xwvhPZ0+0hUkxtKHmfYUzrbz9UTsJlCU03
FO3Cx3IvVlNraEk0EhSmPJvjeMO21SQcd8iT9bXmPFB1t2GC5/+EDxW3gLfAifcj
82zyzj5yMeOBD2MZ6EBQgUAY6aoBxFAaSlgza6F3M3Ikcml5pI9va9maooctks4J
W1XrFF/Jno49CMLRKtRtxC6Kz3TEqhloEaGzsUVidV0c7hI3DueDqbVuvhtL3hVQ
Bu7KJEbyIuHOpaCrnSBbYLha24IFkkOBeSualnUehdH+LN5v1rPwbm5DHt0PgaCC
zXvhZ0ZjmoXDE1gm/UtCQretCHDjcaTHdj9zdbRsxJFjCkOAOzezXasspjDKsuHc
R0Juxz+i/Vslrw8Z1G8AjIunqdwAsT+UhWh6ZKz2xw712nEl3B6/j2PBl807BkCI
0bcjhW1lqDRL8wJjAl7Rtr9c69mzEg/FPVjfo0iS7/2apkUzrHqFERVT5Q5F1Qil
JQ/O6FGITabfzD2AU88M1o6U6VtMk+5hgMLyw4OO8N4Gnzf/Un++SJ8AF5jxU8O1
VcKFObHsIBTTrejcx8tvj4GtjdWn8mal4Gh0RMmiKun/ou6vNNTi5am4XWoKc5Cy
TdNSDdny6FGwFIe61LeKZqOBW/1NM1kUHh57GESA/sNL0aITB1DEZyBxCn4qJs5o
xRW7CS7HZ4pekzcytJbJAMLZgrv0ZFHoyEKsDk1wZ9zFMr99yNT1Ym9SNcYcikoF
DyOYZockU89MMiFXSAmS6unHI7qp/xJDNTPD2dPsNr1O5AbaEGl4ZUcwvdpDUeuD
lzr9umZ5n/qZscCRz5ZNUeoC07+VqcprtSAPHbWxESKofDSHiGdbdlpW/3gZ+ZaJ
oS0f3V0lSKycrYcl3NPXzwJdH6p2Y/8vQVdNhLsRdzox2NoysJVpf5nsI7su1h93
q8rrWV/8GZXVe9d9NoOU3U7NLXMK5nfdegtKPV3mCzAvjFao8NgORP+vlOvfltPw
76WEM2k5EfUXTZZTxpGgd3XBKGkl4ptEnHTx/aXE/zLibRkFWweYlajeDaw4F3nT
ZYqqf0NdVTQyZUQMYOnLE6L1Q0Q2JUi0r6FbheQfoHALYZyj0pw665MSUnHgnHqO
RjX8mL3txMpW7uKjw41bXEChoBaLn6x69epF7EbWcTVINoamdT8eezvG5WPCbQOi
nLPSK+1jE5e1NNikhOZfziE1Lk5MZutRfrW9J8YPmMfVvH/YH4InKODl6rxLhFZF
knREEvZi2b6e7O1x/amGRHbn3jg4Ue5I3GzvztwBdjR2PijOWGEYeG2cCkB5769m
SB8KAkcuMLATKwuXEqxhwhbQQybGUUnMrJx6TBuVJTkSVHG7cMVbQwFFxkqQGRZc
u+SpmWMR69kM1kWhMJRck4SbRGQbctkpWKUTzg/cT3mSFCpM+osyZFdNUCiJFcIh
yFFTt1wla/CcvvACr6BtSU/qe7l9X56vPpFT0/d5ovzM5tICdrNlj8K/oKI6h/gg
0njMFGpYDwQC3h1htx12PvEkFOORocEKSGBZP5hZdjOHiPM/V/1f6sh3ulp9RVGK
hP6dRWuYW9VqsZDn/jTJTLLCGNLZyoEz0ZkhLjVhCSrQV2DH4Tx4UvWCeNOtAEDn
9Np/6QQvR2Z2OnYKxDEx8n0pBYYjX8OJ1QPAdkei9nBUKEQA7rejHOnvzBtWTJPE
X5cIbhaYh7PiiG6s0FtbiYgUIHcPN6LgJ9Rr2DtIHfCNOKQ+WgJzkp72zTNigacy
5VBpeHcIyQFRSSaalXwpDFYF1eJ4pjXSPKDHrfxzomzek3P5ZP+RXswsGv6ALl+X
noxk0A9b1WCuami3LF6Bs1KGsrvkqyiQbuxAzdtOQRShDK7hbb5YvKITTD1u/wkj
x3fntLDdDWRGl4TiZ9Z5XVgGtjeZMJBnZmDPok5AMNL51qXue4VQFh8/xe2fY980
4XtjMLjTxJ9Sr+EXAmn+AuSy0kBXuM4uKWX+VaZZKectTXr1K5X0iCF/sKN+18S+
Jdh1AVbI0L8eLmZ2XXW8dbbi4b9J7ddsp8tELc95KdcwH5ToPuLgFWUsRPxVqglc
ZcMUdFoq5BmLgWSffQdRtuIHcEdZBpETWRBWY0TTcF534tkRVCkv2ypLWdT+22Zo
bG1svWOvCEoH9SYz7mOHKBa8fUZtaujITFmX4jdAZS6Dq+/EbJuTxQfgbIo7E/Ty
zolSrs/yWZXJjTbHh5lJjYgq9iliuGxJcdR4xtD6uj7aJfYJaxbwt1H2BuBqDWEi
ZNNM9DcWO8SCK3S4nad72S2iFHQjiVsUcXQAae1s/DFoIIBgsJw43jGmMj9xl2M3
c5t23whaxFAy0WAnj9nwYU2MKeL30bcRzJ5Br+d2LIDTt6W8EJ1AT8TZxUT6hBnn
+0h8dZ1xMWaPcq2N8kSVnVpeWRZjE5zhrOxEFElI53Y5lpa5c2q2h++UFplXGsGq
akUZJyrxRrzktbvTuxeN8g3B/z5U+nJ3ObiaSHPytiHywpPSRJbpdgdpQM3C8nG8
fOZ7tRJGE8BxoFXp6LaAPtjtPikXPFGW9zeZqx8tFHoTq/7HxhGpZq3rm9qE/uKK
L06d2giSMaDnnhMXsdOl7dvD8nJLHtVPAyeAwwh2GjvCjyYTExqnUeM6Lb+0WIcu
R8m8wSfA6wWQTyqxgGuK/XI02wOMdh6MjiXKU0q0to2hi9mKf83PPeMo3OMYmAkj
ohXnjEbxQjqaaEJ9sUNu12L7iyQb19YBU6YzJaYYszw3FgYSdsFNQnlcozRGe0x4
lPNhaAAVOR84nRuofoOZ9DzLUbAgRZWTFS3iSoR6YbbB9L9+/9hS9+jaeTczBSWr
3K+UkT0Ya5clBJNuMUt5lX+iGHS3+g84JLWTXVZkgGrVRIa9p03MwldUlJ29olgk
6JP7yeGJJ8lH1+aAbekJu6emD+QdNuGVEPgnUAqUz2SY4VS/yQsuUyyPtFYY3/RU
WlDgPf1TUZ6LigOUrk7oI5JHJjCMhPbmn2SLUZ/nSYizuiesRUkuXwbmULRqhT5X
wnXIw/tOzkNebJ8bOfyplo4vXel1Br0dF0nTGiRhwVg0mHZxF/pMiNncFr2Axczk
9lc7a7G2Y35QnVMRaohqgdlUwvSG9GjcxTy3qgvfSYejAiSWQu5z66WJwDXC9CvD
z4z3GOO0kEfIymnbMZ0z5s2g18myZ+B1vTpdgG7jUKtfVfyKdQFNN+G+pLjWHAUN
RINF/Qhv8mhMgMJW+o6/1lQrOtUi4J+t8FNeVWW5hDJfa8t1l+h5/eQZ4R3MQse+
oiq5Tp3zZgLAGqwphAOavz4Hu2GyEPw7Cmbq8sppembtnFac4y7jV86L3PY72/9r
RgqfkxVYSQqt1E1l1Ez/JJelEkzAo2WY6dFc2fbyK6SLifqPkmtTdfrg0tBK/Kn/
QO3gYj3kgjsRnQse0dn/EAzhYG+7gQR7v2XBhIPpCIJiUB5X2jk598P32hOISi7W
EG1CrUgNKL003D6Dt69VryyapUrrlX3Ue/j9W71uAbWxWa74cn2cODyLsBQSV/Xj
6G6qM6y0MTydAZXrjToHRJH+aCRihXoX9RUFJJkI6h0AqnSokKHXjX1/E1zfwwf4
mLId1R22lJVaaZqcwqN4mwHuaZF+ApoKYi9mDg09yvOlCP+9MzmJDNAQE2bOqw9z
H2YLvqz551lSGs6P/s52XXlOyqlUrShIh32i6ZzxxdFwCZCx3VHV/sFAPi3qbCrM
0QlnZEL06dfpj1gb25wnqEBDhOkwb+/CUpjOM2D+/xYq9+s/NLQ+Px9V0fyHqPeL
krEQltC6nqZtzvJ8JISryKBugnwaKZgRg855lyh0VEHszJEoXItKzVokLdXZAbJc
MCrUNZVuhd+CAtVf/S9urSx0E1kAeSt7/bGGaa/8CuUOeJSkWt6VH6ylfxMvPHAW
y3sFxwkzOIqcUYBFocmtdilMjcR7AZxsLfsMBWo33ohD82k4OSAfOqoyyHV3B57z
Sy0+3IUGM+3EtiRupC7RDWwZtHoEeJd/G6SvF7eZ6F2XExHoLEnZbMdhs43gWgtG
bbwfZZ5YBrt9oizUWkq2J4YYFNsshBNlhcqwVTVq9+eAEXKIa2WOphrmFdj8fX+a
HIc9wlkPrzdXRdyhCH8EeBdM/Tvm4u5guqFS/opMYyRmlzp5RdHiDaz/JwuPkDZG
MtoDV9NteLysFe3zZ2nzZrsn7G+z+V+tzs7teqvNB/9YQ9gR81XvMDa/LPiLHfFx
C0qhyPyaeUuMFNkhEQDpALcjus3PZrfgYV90TxV0nMve8qW1SHF0RXy+Rg9fH0pb
v3zigGn1gDmtGihMnhYgrlmY41hly4r49MnbWJi4ziuzGEKHkrITjGTqAGDsROIZ
8NBqTpzGW4ybETLVi6imHu9dmldXMLwm8eP/2qPly+SxzaYPTocviIvvbrdEkIrt
YSu2iqZFDTprZC/BjqVi2rM7OteUWcR2sV8H/M0ZPx0qOfyxsVIaU6ET/y1l5MAv
Qgk/2yEJ5z+zwc/UEPoaGXcQuusJ0rj8z8Fo117OH4Yfgr/oDxMBRi+FTvjF8+zc
TToIJpqUEiYkOTlS8xVLp1/rfYqnGnM/3Ygq5zJaBdvbsIQSHNJhuNZ4HJCY6qwv
YQ40tpJI2zDFEGQg+KnJYP5aFqR07bpEgPpJZUIfydw9hbpwDXwu9P7JN1jsOtFI
FtVj3ChXthNUdXwq083elih3Kt9Jsv2Gmk2yMxysq8IVn2VEqXOgz4oXDsGZYrhS
KPt9H4p+IRnYdNZ0y7WFKvxCBn210MSDno8jR9wdd/eysgU3imxJ+NRZIaPXaQGf
U0bWoyLVmdsGwOJb7NgKJZOAt0/LOdX517SvxZ9DSt6toR2LD8oL2UQ62ayUm4ts
AgPu6M8BjXShW9QCYz823SmCigZTKbyJlpm0g3PvAS9PxdQgqKax1lsaKqcumMX6
CP6ITqC4XF6D26ftucqRdfaZk2rUSoF0QfjErVx4KqekfcTSYTcBW060c8xBvprn
fFGc3tq4ZbH4qJW57sJLElzenn4ik8+ixr8JXV4thtPIoSGza9r5QUOdsha0+D50
Vth9to2jQd2TPEw9YMrDyeGojOVp188ofc84GfDImabF0a0/4bp/iiZDPzlpzVl7
3GTcIRGvw2sH2EI4t9j5sFIpANS+8v15v8tZgaih0+kfRQHjHTuSSuC2LhLp53G9
NYB+Tpuak4JlNlDJmKxfi0ooxviSfVZs9beoa1e7vBQwJhze/2qCdBTsVz6Nayqw
2uGBA40SqkoX5uGVtoWDOOk7Sic40AWNt4AsrBaPJfvuY39jxM/UpblDD7w8CO5Z
JUM4injj/WhDO0KIqdDGkjtW3AaOCq4oT4iI0MTurnHUuUHKlOIKQefo2EWwoR7M
GiFuY8U/em8ij2RMz2ZtWqbxagyRaJvHX9n8uW+/cQOYdjhD+OHBaR1MvzHJZrKl
s9PXy65o4q816WMWv8i+sf/Ryg7ldeiyEk8SwRGCoxRKYPJTsWWa7uMhh+PDVgXU
RGvysdI8WhwkpFx55FIHB0qTYYzx4rTzAX61wT83zF6GOW3Sq5Ite3KLEvWXVJow
KPz8vXqVEY6MtbL+k4/9vtL3cG2MLFzBs1jduRVbS7H9/bsGONsu0PIOR09Qzedk
U4yPLIiTi2IsTO32RqQc5fMjeRElnNkbHCCkJBIh3NPzIWfGWr56NY+IzV+w+HN6
I/fT7ETvHhfKN5OXRLTI3OG208389FiCfO3YpU0IeCNKe2gOewf9F4HqJKoAo95m
sIFnRrZEh7mpi3Y9X8YPAPDx4d4aHb64/N8CzTAcqkmo7WsdxLhCZb4TCJjsyKhD
X2BWS7yp/oTDNgFwmH31jXIsc+z7yK2zGDCqRYPjMXQrASpEZ3AVF8RCPSi4Y0WZ
IaJA9G9cVV3KJlkLdxzJe/+vsCwTmDbTiYi8tlALdtEn8ai/kdLCypgzz6U/3TrZ
FwKegBnNtye4koDWkCQZCRi81AueZQRhMr3ZbUSrtqP2zzu+nYwVR8te2KwlJQA4
PeYBmepOTzk7H1XZ009Y3xnWBaPTx7EtPJpNPZ+jt9bjl9weMTgi+mBx9D/XVino
SSTjs/z/OCJT0vEo9Ko5vn7AoPHNXrGVtv8ytBw8KEfZKNK9G5ZgWPfVAADDXLco
Czoz7rqcp3hIZ4e7/tHipnxe9FLPdKG2VaO3R3Xph5s+3L89MaowWH23EnVBnB2r
DNSeuFEIbt2AFZTQUrNnJeOMrEf7L/lp8LQePl6wquAicsKLGSGHV2GA/6fvZLsp
hnYtVhPxX7c721ATP9KT/baVgxm+QRFy8RDiUBRQnx4umkBP9Jn9+6ZUFMKNVvxE
0xjd//fYjIS9mDBUhsR9n2szy04zBWKTNteU0k7TOWwL9Zu3DpXpEnjPnYLOEYky
jAcc6mawM48UZSuNrfgc3pbvZsTTe/3Uf7Pj/NInmj3be+X4QZbg77UcQXyc/t9z
piyFn1u19g6sI0IPtreXSbUckq5yFvlrmkVPjGiTBSia5IkqD+Wk5Nt4SxYvgJEl
agPWy7084KeI1RsHud5RM1+Sd24I++AG1sZ/KZiY6lgJaEbU3noLa0DX/Sf8GXxx
P5680L+DKD8sdKG1iN/4M/8C/2UjvMV27CkfB9USPVkri/GPjjgW1jUe0QYkQ3EZ
dMo7CuI1rOq0h4u9jq2wpYKVU+wLsqCcNwbzpIC3tpRmr7yeZc1fpuqtEmOM6g6Q
x1bcJc3FspdeDaEnj2CHcf8OXgb6A3fpXbzZG3YrZ6jKzkd9nGBb6ZwT/tFSBq9O
kPthHznTEkIlNtqdx1SYuQuDNFJhxDxAOXb4qz43mV7yOZ0lIL66uyQQPaHXuu7V
DdlcXrsGi1NTLZRmZpR82CwJuumS40D4J7oipohyTRe5mWIta2H/3WeUzvnk0zBp
GL+fvJHwuRr6RmBwtAHDYi37klw8ppIF35w7X3t8S2mTHWoSDkYPohrdW4SXCqLZ
q2SqbGoSb+Vd7IFto55kGDlGFsa6yXrl9bI7k/hUBf1Ic6GV0B75RPgiT7I5sI+Y
kLOefNWCDxGc8AZ3R2lr/vx4KQQHgZmDuLZd+ZRk2C7iN9q5j/vh1zhDVVLzCxxw
7e+94zDgKwj5u0d8PLzIhUTjjF/Exfn1x7JRsS6UXZFZeKjnzdS25tg19HgQlvUH
oRMRAYe94ZG6PwiKD+Ik3eLiJlFR4NP6gqAs+rS+i55WNa+2MY840DApS/XOJ990
aug73UhYJrA0QgGGlwavj/Ts2ifAgWH0ETJL6F5GOyJVLZYgO/b6G31Rblg1NIGP
PrL2+quqaRU1EE39OnMRCQYsC1JXJ0I9bRMAbf73d9iCOap2hrwijQotjDfCCcXl
qEiIExns9n/UFoPiaxSaK4kCQs/YPC2lMCtFUVbLBjET2TqoaWCMsxgKYO0gSGXy
GMGPqFHY3GPmiLpsdXMkTSelaLr4j1SEFNwTh6WE74hrixw1k/yfyNIEGhduvex5
Ip/UFk4hP5fcrkymfv19mUe3UEttQk7ARkjG/lTR6gXzed1zpEBQ54PqVjqULScE
BjlGR/FC/k2odKK27azFB+hsWgQKG1hmGOv6Z+ZXhy70XYNQtusC+kifyweP5WXN
WClldNP1eYbGhev5lGZogwVMmpcITYKrdEdXJ7te+AL1b9bISTFEU88GLqH/YWIQ
LiHKCvvikPQrWX7tt9U9TcLy56EtqEo5KWyGdMfwezCfUzDdmEeNjYpCHmuTV1T5
BqO2FMb+a1+FeLubCiFe0BKEFmVLRtEF04Gtrga6OH1ItQAyiMeCtjT8fyrpGwA6
UQqjQa6ENk3UsOnwD+j7ZpwxhBSKNjeERWY9aJWZ28QXfxjXdZa1554w9rRHNipR
Gs9GYW1bk5IwvkYCjMdvSGdnkyPXMixOdVIJjkMn6awlPgAk0pDYubDbH/QXaPof
lAfsN24FzG9+8KrXCaU24Dtm7fQLxDaxAfTvqNVCELi7wM6NV9DL9HEerCbuiLRZ
I2sYlw+BJAgIyF6HxkqYGB0lI+5jmv5D+hhn08wsfFIHZHrhssljXItXOAqwm6iW
6EeQBB3RdTQNTJ0FhqFdlZcEltsJzaQFMHmUviaL7LeusYrdx3dlnPqT62nQUQHb
fvtRHub+XhwnMh9+v/sxpiq5HOhiyhTG8k9of7ourcCUsQQtBJ9MA/I4c9LaWWxf
JLsuCvgeLG8doG7KwEUy80SqCPyuwwkVzkXWy0sQzIhKrmtUev0S7jwMrdZVO09S
QKGbVF5VSvs4xlhbgNLlJIdspn1YFxqZ+4TaKF0CPVJLJ3w2aY9McvjC88vEYJ6A
cS6jaOUpLD9t4sa9kU1moNAqS3eJRKe2aIymjxERXDQ2N9HA8Vvuey7D4EFfu7wK
9KIad0cxzJwKok/kWLDUmmoMiaBUFR7UenXNTjPAi30II1rS+XA2f4vFwNL2l21y
00JlncXK96wsvh1c3PK3SKVaCVfSrqiCdxsStjunz1SrTAUzUJyCFIdPyGLPr4MY
Hycv092EqxU14ATXChQ6PzjZqaTXjLgxCJKSBbQdcLXDo0WoGVcX8+IMFNfopZB3
QXOnOkxFbVq9gUuEXmadjcHT4JHE0v2pw/Xd4ZmAzww24N7NtcQX+Abwst4ZLU+O
og2bGEWUp2Haju0EI5e09B58IwRZAYGhnrrEmLbH9cMyB8Hora2860JIAOX06GDK
7+c7VLXerQ50DMzGVTHLnCr2UIXD9M8kSmkdr7SkdTejQ7264H65funXWr0usLHh
mmy/MSp+3W3nnZMo5slIjVE02O3swkbvtjSV18NBmAFTB6v3XpVmnwObVQ+cdsQw
yFjIWWQ9aUiYovG4bKPhIKxybWLqgQ4ycFmfHLkSbj1QMy9Ry8go0tS//afGRNTv
ZAXgf7UvJCV0GxnX+SYJziXrsANfdFDH7+XhOMk5m9T6s/VTUintb6WKDRHG6KID
ufNv/GEEWTr2SE9QsKB8Bhl7HCLmOWXr2GhcanN5fYOTjluIWV5Qbu416ZStJqDQ
a9tkV28sV+HPfu/FK6Ap9yWP39UHznOblh+2zj3NJ2LaA1yn1NvCIBjsGkredWTy
MqnRXCHgc9qrD2n/kQivY8bTpYRoZ6HyUNFQ/D5EtnmHIEztYg0cKWfnHl6nrK2T
0HklrHbM53a42GEbhQkrn+BPnHP5M0lxCNvTFcVPHgYUBibOg+YPtgX5THLwDnkh
jHhP0hbJCzrgpvqbQjtQ+jzXZDDBBA+ZgtiP19g8tY9KVn0heIn0rpEf0kEtpkRt
smltRRoGkDBCH55ksReSC5A9a+AllQC0bLrTi1JS/RL80lb6OJ5Oa7Y8VU6ANMvh
n6Kw+vgPiM9lx6vkY2E87lPU7iCEYWKPMb82GsCVYZcVPj5zmQcQrs4SnE4HD96N
aJTHYpRgqHidpF35TlmPXdBlyvVao2o9zlSFED0gpZQxkNEbKSoosa4ytsXsmttO
crLpLdJZsxgxStOWrhjf7fydUbvI0iYv/xDAHhDtOdBrmASs1vQGOwgfL5Rkd+mY
osx76LKQXQIVPfpmOo1+OBBE1iyaeYWZvGMSnn7y7BKzkU/u+DPiheJuoZoggc4a
gddGbRa/3GxY4ucbE3Zi8vFdVw9gG1W60XJnFkv9CCcVE1XDMmJYcaqOg2zyr5+T
zIHOWDgrwFE4tlP2/pi4jaZD6xlv1JpJrLuuXZibg6qX0XOsTqNPSSih4Zi2agDX
2a7E/Me10tpUqgrS1PSp+3Q1+yAT4O5Ls2fV2DAhBn8gCdf1dfTIpFdqou4HthnA
sqtRdn654Olba4/k8Vm0uiLUDqNW0HqHZEC3pnS+U2brEvW3RthNQBt/F5B8HSJ6
PSn8J1M0Nx5zmkoZfjNgvvO4Lpy1kz3nmmlpJNgSOD2SWDfLGokyxFsioRVI639J
AkcIraZsQ8iCJojU413skixCfcPtZvwI8nIIAcXq4iM5A7Ua3FOcV0F/prWNLRc3
oc7KJUTUZjvVQqv8e1x9sS+VpUa4qBGdRGXR6pGGX3iTBS07+l6CAxH5/DYqgM0t
Y1NRYQSL5X6AnEqNKSSeYT22z8yz2kmvRcHCT6dCyS+M5sCedew3WWV6+PEqgAcT
lVKmBr9scwZt6Yjkc4i8sFVzhskcN+OZ1teCa5sD1LHfp6rRWuG2AmSV49Ye+BoB
hz8WVBuikld6z5cZx2IAJkoGcz6XT52/z56FWJlKmBfgVKxfOXtB9VR/40UmfHCH
PQi89ooZRoRJA0pL3lnv8nSDipJdGApIcky0rniwKNjS+3YKtGC6w+wAkz4XW2hN
zIRwfDHvE8ERHpWioeBIIrmUn/rR0L0SfsDNu3aHhBBBeAi/ugrgWWkfEcQU9Ycd
GQoem/yZupfob77p/bkizAeBXcjMb4E5C8EOzgbaJRhjx54je02nIbyV9vTRd7Mt
4f31Z/qCuCCLfr2dIiCACOj8lNSZsOnwoprUapISuiUl8Fb7x40LRFT87WYPgMW4
/Tm/QtrmLrj7nW5Lpe3IK0oPUUyphXMwX3dI/QmRo8uzr0ZWEnEFAX/1INEjeUQb
tt6tImMbBWxV/o9xzKz0IzKm4TgjWVVluoAHWsSwFby2TyKQpB/PG4tWF+skzi+z
CZcHDTkEDpT1v32XS6adccMMhml0Eg66PheWc8abnLWOYsGBB793hHLPbTS7Iypj
FeFDXv5OzrwX62er0eMhPsU4yyr3I9a6OW3IbmjrL9DWINQrHkwQVEmohdH9eiIz
bkGJtICPhgLsplTcT5rtg0dbeduafDFrdjBRRLCarH3pCFnO52iyTXYa0CA5414/
58xL7S5J3agf38zxo+x130R5M8df0l2MHHgo4xEotiHzUPmhfrrEkWlE2R4qmbVk
hLpTr4qWhGso114Yxm6lEyY9pqqnRWuMhSldhDmw6E8GGN7aRjcHr2tdc12cEklC
XcqTPc1RkA7FQZyRRyFi2vWNcXMLjB9qbYODbD9f8+EFVBZ4S3XWhaP0K2yeTDDc
Og3rnaCKzFOcoJGxm2uI6r6jI5bqefiv4dFtuHXn0bEXaXLYf0UPajJu5UG4aVG+
YGQRLmLdeZldsiptlZVCnvyTOBIKDz+2exCYS+zfvdYkX9SGGHwwkOXiUdcH6/7J
YiMgtgo4gLZIgES8mt2Acb89lW41BmpCcezafsu/hGjfIw0eOICmHy1rj0aIP4/z
bmGPO/b3FjWM0oKzyKQLSBbbBHEFC0xsWtrOgXF53xsyuRMmxAiTSZ7rGNAFQD1T
KhEuYqd0S9NRUaEbJk9NoEKL24HuvBGzYekLEUdKVBhCVugQF90Q96IJaAhH5ZtI
lN0cHOmktntWh3n0uSdrJrwGxwXLyQoFJhpQdSmY5c5pxwF3f43vrzBkf1q18HRp
sa9/StthpkN8/kzxrBdkUfZ1BQ7090g34qNqE98D74Elsoev4t+wB1snBu0kffLs
QuEwVutypFuIV2qSdM/3XG3Zwzs2VCVJTpQ2mL4T1AhT4MDFqVP1zEUp1CXHFDyB
vuA4lDHiajdTVGxcmqglNM9DW3sH18le/cFCDmKNqPA4RzwQaFDMM8w0weillBv3
Ikgcto2d521MWavRXwx55mSDsqf0wfia20KNcIcONFfatUgWJo7p0HMdCk7IpwoB
sw/YQpqimNu0BAeAzXsw4HUXyWlv+23usc9rNpzJy4ReQF/zJ2EXv+d6V3b/Zrk8
NMhcruw/h8JIf29B1hog9tiTdG1qM6e3cseIyPrO2otYz01RQ4FZmpLaMT70BpKM
B9tonhqGe6hu6vM7SSl20fDxXW1SSJsxZv5G4ulwg64Q73sUOR9KRxCrbVjtb/Jc
xOC5W4GNnQZAvsyv0l27ND8/GCT2Nf5vURVhs7hZspMVsnGwZHJ2gHTWTpDIr6E+
iRb+4qLA2wFlbHuXJiqbzDeSaVu2eQQ9mBuBPzhs8S+K5PtVtGIhe6FZLPlP+SN5
gWSiNeohIjo9BvK0nO/Vy9ZSOnMlHQylr/g7Yp41r6p4iwCRPSNMPx85CH0AfdNv
4aaiX1CDW2Ig92eJMaKoGDQm3ZwbDzucTfZIABMpDHitsTs+BlPMppG1cvrXvjES
02bvxmzZ2l9TyOlMDwbFmPomAXCgilcbl13nLWxYLKP88eHmDtEcaZTakke7VxPe
7EBvSrULU910zxXjhkhhUZXKc27xooBbZWijf4Hk9LX0uL3Mj8QuL9nvf8oH6RtZ
tPDERQkC3j7XwEr5Mhz6G4QCCn1z5uVnwx45Wzrmj8lZLGT09DaNXnHcBCEZnWFF
NfH3q47Ub5JRV5Tnm70bMhV09PEUm13tLF4snTGGlxKstFRQz/fq1d2R5EvWsk5m
OkSyh01f1uzBNBCyUTQCmu64k/13RU4F137rORZpOReJLTWjotEtvctZoOKWSYol
FJU0kgqrvMpl+OWtlTMmCTzpSa+5wwDjUOiie1giYo00NyhHa6BcVt0QfXex1f6d
SqTUHSamRJjuVaHN+M7m79ixnKCG2u0mZprksnEujWKCg9duWGoXRaf1rTQ30ZsQ
Wwx9BHa2qtIbRZE324LwNMS/OSzCg4rS8zcOu0n4QrREnsXHG0feE/B5MaAIVd93
v4LfbcbeM+6ItWxaH5EHJz3lLwO96+T7nqpi6auZQfdnzYfTLL4VY7JLjoUi98C7
8jQsd3LBIalSnRAjLqSLjufhNCQ8oMRHgQHLwjhbbIiTs55Plhb44v3Gb+Ua3ZaU
Dj8VidsRQyzPL3IrUHnWdDr++YelBHni0Dk1hsKjkXNZ/5Vb0ZQpGVlZlDS67O5Z
3AOJo5ezw4jBn9++i/jdV3dWvHC4oyCiZRqbrie4b8WxB07kk0iHbOeuZ8oiZue0
WDWluU+oRXEtU3TUApHuu/+32HgH3mugIp9PcJggkbR8Jy9/+E7Nh2ttWEl3o8L5
dIbKUSUiANRXbhdHDZNGGrb1EprIpp0lMyJQOxty4GzcohEDgVGo65hrWCoNVXqG
IBjkviweG3hmJceOgX40Tr5mRY8JHRhtjSIq7Xx914AbpUMliOwkU7ETEwUyYGd5
u7itZJpXsXQEX0qggrftoJs/GFjJNC04UJEorizUrPlXHWPheuukAYwGIgWlJegC
ws/DAv2D1VbUgIGqkEHMeKrw+7kQZZ0fjLPdvnZdtQjUCNFULu1YBbBEUQ8OzuQL
397FIkHH9jrb0/q5SeWTT0ijsOKLU2XJw7+wJSISN0/GxVO2IxNT61Kdy3dyrPUG
AolRLdVn+/Ptq7aGQMxtRu71vj4RuAoYPwDQ1FSKT14ST5UhQFbBxCQp9tOVH98W
kzlqXqgWJMsLXNJu4I2oelU+eA4aJgZ/k4ITg3yp4ff6XRrJJKc5MF0FPNkskAhI
kEpHQmu0lDbsTjscsHHITy4B2NezOdeWGixUEl9QqD17HtatsGDEGFlZSU5oiUT2
gQKF3vJdl9cVq8fY7cLEtJQtsG14Vd2gamsD4ZKfWXW8XqDUp0W4SMZMxzXi00Qe
KOcXFWz0D8whqIHLFhnqd+KQnM7k1zPvrK1kWX3AHH/mtUes3mvTkQslGjImcSmo
YNFVpMS3y5m9TW3kMtSqQgT1C74Dt/r75Fw5ZhafaRUXffwfn811Y8d32qNKs1jJ
iVvGjknYIa09aW/fkavYyFxeYwHNvifsyuFO1DqKVTA0WXZLGTaI6YDqE63immSS
TYsUcKsN931Bz5r+LpzeQNIYuf9wwzCKJD6fUuVpPO7JVstUrbq2bJd6WqXQpZtI
I1IPLw8vc/st6GHKMod0YXQMCX8OywzrwYY/I1aVLWav0WRipaXO6qqY9013d3uM
0by5PGt/BGTvY/qx6kSrYs8fyCbKV1nX9uP3s5UdA6BunKRfxYwrL2aHhNQogInN
KPKBT5UsI6PuB3N4lwIlkX3EehUruAiZP90l0Xfjhgc1GaGLKfcgO9ADK9N4Cl+m
HZwg7EeHQYCkK39ginmFE5UVRTVgUK13U5Z0fFxd2PsTaPYk4a17wVQV54/Vaw6Q
3CK9L2KQl0vVSjh30p31xIa69tWQSCWpTZuldognNczyaLntktK42kenlr22rMHg
ZslX+4JVg7QLAZd7yysMJK1RjrwxzC+moIlg8K4LnWjazF9yLOjVeXq2HlfslBwc
fHxaWfcd/2ZqaRkVsOtTcFG+y/s4sI4V00FEpyiPpMwYxtZD2xQof2mpeIf/tvrf
ma1sS9Oz5zN2sO5kZh0jx1j6k7FrHRoxNfbMDPaN18yuRp5rXS2zR+2r3NiIPuBl
DhQmqaD8mHg1euK6KM2D+aYsGvg+0qO18nVTFd2302t3uI9q+ldOpwaOie3k0+Dk
shcHcxPVjRy3JMqsTz9+kqpSKyf2LKxKClrJxSHA5HY9hDjnBkYI9z0j1J+nOYe/
bYT1ShRglxpf6HHYA7UJYhzb+C8ewbzt2fFzbofJqNlZd4R5BKLxyA9hmzo//Rl4
1bdzeQxQKMi+AV7dA/aYkfMB4JHc5KHJrmd1cCcY/YBWzEaNq0Y28H/vzEq2FHct
g+3BAwPx3iCGPiCoIgbR3l3KzPhVZSLsauxY2ZerF+DncaXX+2EJroUDRbtMg7WQ
X3yr/LCopXVPUJImrzy4ax/NEzeVSFgm9FC2Y1QU4rlT1zu1eVTOj5nQ7kduDNfT
Hx+kMjBxvsrOEPsk15LIewNkpPCXCzeUOedwLsljVhPnSIejagyJOfxbe8zNhj5R
oycvzJ3q8DybU8CH4dqAdC4Mce6mPUSSV7JDKVD17nCsZ+dQWj/f7vY6ddU8a1M6
U4gG1x1sWa9oe56EPf+xuMyWC4JPc2ks/Eby2OIitbhGvXtDCXuq5Eysb2o7g+Iy
xU5NURuu9Ampsd79/KyxJdHpNr5/CCggxZrfWADF2ry12l+5BacijyzhRlJsI9PB
u+WBLUNaY5ItgZxXsoFjQh5DyO0MZbhyXrQKJNXrCq3zxkXzuueVTV1QMcMN9iu4
3xRMHuXit1CK7rxSQKRXcnl+ZByGI26B5tBRmWa39yJdTqEvD+rpzFLprnZpoLTf
c0S7/FZRZTnxjxpMwT0uSUV0H3+2pSaUJaaaBgRzb9hvD7d09bbIwdHCxUrEzhJE
OKnCCIleLOtS6kXgwFFtNQFed50n58I10ek7sZlMK1g5ieVfpt/tbCroWZ5/3ArK
nwWMlXn1qUg3SSqo2Y54qjXwBPGv8sHITvx1bLDi0iIzNawJMxfjUTbYYOsmZWOR
3/BWm5hnq4DW7i/Vt3X4ayMQZYnXAgbPSX18Jpxh2J7iWP2XGapoTzcoMTpUaXX2
jb7U6DJUHiuei5td6bhXButGmtNqJeY0noA/p8iWTrxbgEf+ourHW6CwCBZ0wieJ
12NmKfXe3Z4Hk0qA/7y3vIdbw5m/t8gqYKdyn4gaEUThdba0WpKG9XO+lHfqgXd+
YgbLlnF8784/fynOD8tR710MwGn45ZErHJ8p1371PGNkwx6g43tDHOee8xqXQFqL
AntLFxj2+eOMAbIWH3tw7ggrVUJ0flDbfBSsUVYExmDb/n8+yD+BWsr5yJvKQEPT
3gER98slmsMpy2QHsFRXSpEPAsBwDogNUri3yJOkoil5LPi/U9+dnmVHNkOwX9r4
50CPiL48dySf77sOnnwrSpE5GFKUb9GCi6PyfUmFh+Ns9DIBwmeZMMWIrfbnp87W
zuNNG+gmXBHlBs29l25NfUM6sle0cOUTUUzjykHcI6Co6IVHTBsmwBsNU0rvzq3I
8udBsk8mK8UyYVxbhymbCTV2IWxAHDvGG5O8HJiTRLw+fjPHHkZwEhYPH7qBgrxg
v4prHQY2WgCdrQVe51wNwkk9gtCD0DQIxXm95tadeOBe7Ln6/crw9BkU42clnMxH
GVR67lIEhplOP8zSI5QHsLLL+arr1/5Mtcuz9aKGYVpaoH8/Z784M5Qm0Ohr5Suo
DZgSC/00Pqgsm7UXrzOEi/fao6U/Yu6umxBrCfSvCu9sEBHPOdwyIknROBOhJYNw
893+3CAPcDaFlWDtiyyrptVvQwqbhplcout9V9IQCzQQkYsk092v1G+KeTFoMzKE
zvw6LWvGMoE2nRNW07fZxIjdrFCg0EGQhlz6fSeYzmyGphRLovavuPI6qUxR3i81
h+CptXAI6SLvZ+lS/XJLaRmRZkEcwPuiRKl1//jTgKqyfO/isadzSpjYM7i4cRAu
l2dz2BayvMajg74mMLjOy7nn+FLK6fyZE0CW31qD3PkbjIlyfF6pcj437QsRCcgt
SNayNa1ZeCG910IBBHjim5EqSyWUJa6OVzLu3XiHIllW7WLE79nz7ZeYdqt4n7y3
0EtSMvLScgNjei5MAXVkivrGF7l+Uwb+ETMWC40gylUX2obrpBtpHkN4y2att/IU
MlQrhsDzUEsIw5eyZ63JoH8+3+4Msl9MHaKVQsMVWXsAQxjZV6DTR8+wpJHcjSll
jsedM7URDHlOGHV5Ruh1/IhjHt8FVBo8ct/r8XdbEGKsJEo+sUnCvDZOvtOUItzF
MfCX6f0HCN/pqQmTCSohjr596zML3Y0kQuWJdxQAh6+1OfOghtE6xjNvWgwh6C26
ldVdZ3xfWA90QlAusIA3NbzLOndxberzKpbhdFw1sEr1j3cEoloSjSP03nmG/gj1
+fGZ6GHlkMif96FFvFgO6qkwCVtjIjArEOGW0NPXQRtxDmN21H+iDpuM0QYTib0E
k/CL6x14gJkgAnKElNM50pZlKd6+LxO9wOLaqKjzNFZBND3HuNLfjGwlrXmr7rGT
ivBwDeqYaiDUPmyuy3cDzS+qvFMqsJd0GrNNHArbu73LCcnHfaA8kh+lXjUHCH5H
+trIAPS+FjWzQLwBNOL0GLyEQH6uPuiWAs3It+PgbFULGBpED171SEnYdTFDZz8A
sLqLQkdgcNQefyrzoEekkkcnkOuezO5sLXAuOJ5lex4NJfKr9dxO+yBuHLfVGqyE
Cxgzi3Bs0DuIieIctTXGk1uUUjhg1vAzAUHR62pQBrMO9taV6mAWm/IYyU5HZO7I
dIlL3ccXtTCMOc1h9PDtBaDIIRdEoCRjPdHW8xiJd+0xl+4QzwF20ivcxwVsqI0v
DePib/Nz/rh2Ei1YSWc2VP2HROGJobILGWZeki6OCcsJAZN5oEZqlWWgpTAw00gR
vrRR4+LitzCHwEWBqgZGOrcZQQpdMJJNK/xOIJPl2c9ODBEYt3xo2ygKtKbwURhN
8Q6q+kQfMwLGfW97w2BvqGLDeOAlxMgxnk0wOLphcWLdgoirkMxhyXftogQdsiZO
Q3Inh8tEp57uyXZowIPDYeOu0z5lu8n3geJReQMEDP4tCb80Y1+tLbrccXAWDf9T
TxhZmg1zTUEHSpkSXIVVNtkhaQbCHZ7NETJr75Wd4yMCtAe7GP8FBROeRaFIttf9
XoTCJdje5NNdHsVREq9olE7afuNFKlhMqlF2azUTK7mtdhk/6lCZdQ/9sCBU0Daf
sa5qiSTLFVqjPuqMwKFIHOG+ulGb8Bbxb5YicdgXy1lSabaqvZR0/MObSVOIEXSq
Kukq4UOU1FDG0xII2cDbXnRR6ldr9KSzItWlpRQJjRiDP6wPfU8z9itiodhujNjb
MimOPdw1s0XeI8vxLZtdU4ZnOQANDpaQZLSybbLmyemJRQXFVQFn3ditR98oG7+p
K3nH2QzVUZ4bhz9HB0erHO6F1ABZRCcFKKbidpuB4rmCJQSpFaAd3XCawdqfje2o
l3LBmc0FeFMnsDoAI9C/gSj+U7bCtMXXjJMWpk6DKuYDliuFHzrRjlwCviN1k6CG
1M6cS4Z74hUaSDNU7fwe6FXNpdm1TAWM4POX7vN+MFATojk7MARD6YGfspOblffk
bjOlykWsZ7b8//ZBDgCgXgxTyB2G/pQhK0z54pQWzBg2mh2p0u+vuzEB8PXaydRU
4DIwUiAuYflT3d+vFBLoPvXc9MgsnYX2xdqj5gscrF5TE0pw0WAfokwamUdCXa0i
piZr3/bcgYvHWdVWYefZcmxnvByyQYbUBWBTxEkgqHn/QRdbb/82YybTzO/+k+lE
YcGomxP3A/BChMXPKNgypXNFdZSyMELSlkcyLzrFZVW8KGUlGYQs+dLWyOWyfeDj
jDS4+21ayHIVfizPuJierR78w2i2Z67lSMZmo6lfaALoGgMqFGkWbL+YLKIovF5g
tYR3KHs3lTdz0zRZioDVxFpqmi0XTaZd4TQars62sz23VMM0Fv1FQCStKWDUk+vw
VScww271/mihUzhvZ0TR/jfYeC5u3tV6j9fa6FyaCVirlUm45TnP+r8lPUn38yea
OiI3V0B9rnvEjtxjyi8ht7JrgAU4sVlTAxb4mWyKWFBMGJWwVIR119lbBhlgxWay
dlaaeU0kzAb6/XVJwin4GbqmF1HxWg4p8JK12q2uW84nSLwkhL0tkdWK1SXZpnqZ
8Z9WwsngutEKtfFFNbRmK9yvW6XaRQy9iDncnyF/CrIwWWhKPMQWLrlZVBzUNFNB
qEgueskCwQTUR3/oWPr05c+3VnjSPPqmxLs0kEbqwdiNgjg3ONB11FJu6f9nGUAa
+FFwC5/F+YbPM7bKorWi6ESViYeNIJyI/c5vXjiu2FADRZ/cFPq/uAUAGYTAMr0M
SQj0SQf+OqYBgbZFiBUI6hlDHeHfuUHP5geyUILulZVUOBwFi1/8xcWs6+dgawAv
cWVb0kD1iP6Acjqjs2qH5Q5YlI6ZfeuzaUss6RQ9vcDrLLYcj8dRhNT6hljUZt3x
sJOE99LWxwZ/wMPkO+RxyleCJSDsrD+XjSAugklYFGKupZtJ8iV1+b4yaYuqvT6C
4un3pkvhlVibBZDU+e97L4PtEFxRo8RsGxZPUofIKbhKnRdw+Pu/D8ivbcKGsh6K
LwYlB5I+2X7OmLBiTudNZa7GJC7ZLm8KqzpJK7A8VfLzF860x2ApTcbwHe1Y4Vtq
8td3EZaRybhk5Sk9C/p1+RdeCzqcASe3k5vke6xyVjaaSJZ0Qgf5ZtvwzorUU3E1
3x1O8AQx2Z0IlIW85r5yBu9y/8hzXBQ8jViOuFrgbh3/UOpxCAokbRAzntPYOYaV
w6f5XiKuFoVWpNGn3aNk/atG+ppChb5/quLChv3YkHoBdHoP0ccnhLc08TRzYHZz
LdlExz8GflIbf7/SdgzNn4orttVemj0pO7pDC2R3/l1QYD6BGorsI+pU6WWnnARl
qGp4j/bCrjR6tEDUDB+Oj9o7GgEoaaYg2NGoSEcgt7juBHSgpz9udliWLTwLJZyY
H8s+qUS6h5Fv23hg92IrdQTumyMRq4ZIskKA1uxcdrHa3lt6yvv/WC4w9vMb0u3G
dNBZFEcrcvdcaOT2YDS6W3J0GXiHhLDHn5Z1kkWdXt3WUN2UGcuvUpM9UGDtVTRM
W+B0OmO2y0o0EMo2BfvwEVlIhTuTsYBCqEVZefZek4eA+2H7gYHVXoDD1JBEDfxc
fUZVwcmGjNS7QMZjscG9I2R0K+FP1jnMLh3N8mIwGZkFN/5dWxqpQrp2IP+dwXwn
Fl35UvE/7t3xPdb3mHwhDexPyf0Ned/WmnLJ4XXp1T0LB+I13UUgeStK68Gy8pjq
hxKYK3VGHBNCUJy71OGRAiEz3J4K+JaanEtTgA6SEye88iNS9c3ljUtfDYmAZQKD
i+hNDwYTOeNWMDkAFlX0ZDb4JkN9M7vGB7c3qCkHtyY7XNFQNFGW4EU9ggzOfZ96
irdFGRpWO4/Gw0QiMlT9MqTr1CBC9vIbK9OBxB6zxa9wbwyV8LjGNfdNTpTU6jP0
hfXlkjDRAVAzT3nAxdJtJ8Do0Cu34QNMFMoWiL9RSpOmThWpnvTFQv73TWMgf320
8vAIO4inL5GHzeyRLBs5myeYyKeMM7iE8vlnxbQIXMnjBeA2RmrImvzIaRRiTIzK
w/PyaNAqwi5esBzYrh2kKevzaTpIFZCkuM2P3vhAit8OB+B4B8VdKe6V/Vp6FOP/
yVPc71i0w0jeCIIHwQ2gH+ATyZdV7n9Icd6vX4cq0cCH9bxsguuqlpytpnJymk+u
iWnlRI3UwEpBLT/QrI3FohkVkjJmQ7P0KeZWxnxKzpuL5dyEFW5JJqGHDsbuFcFs
HtZdeQbRvIqbQ3hu8yK9TEwsRtPJRuHFHozQIZuKxqA8scu14rVF6Cm4nyEicpQL
qG/N15T6Blvf2ioFHKq2wvccm1Llzd27vr/EVtuqTcQGVycChEe5d6RAzFH6ZjiD
PPG6jEzWBMhfGLYVnYs5GCGztl7pUdeyf9q/18hZ8O6OEVtPruk3emW06r8Z7weK
iJqfJEukwZXQpyt6PNNGky3OZeveWruytvFIxQYY4PJXjzeQ8U5l3hXcuOzj8ICK
KOzIrhbBPzabSORJd5I7mJUvSNBgoDbheiqB8B06T7L4dSRpO7Byibv4BxnCfSEl
Aj4Qz1DRDV0KDzIwCE1q53YYW7CmPrO5zsOKZOrOdZCi1U4QkPVEOWVaVUpmESFt
KIFRbMIAjT3yHD4JrY3F7lgtPpyF5ndp3zWa5MzHMCz1TbWZw3+y+0Xsni8giIR6
59+E+IlgNyiWNXgkGp39JRKwqHPiGhxEYONIgHuNGjsecWjYXnXCNWvyf4KkEB4O
m/QZkau3WKmmkxOtP1ap9/z8IkQ2Fwc2bWFigyjfVt+dI+hdxWgc/Ukd1NBVFEz6
0wuWfT1g70XT9TBvhcDTAdqjnAi6zLKylSTlx2YhqP5jm9MspNPxpNH3aAmGAH+/
G4cs+J9g7W93APcRSdDuE/iwtiH7mNVJy2RyC4xUl6u0Pt9TC9DGoINzvJJLeUe/
cUx+2AMhq9n2j6Co9nXC6lJ6QjJhRL+hR9ee0LT2Xk0wsQGS5LHoTjmfjKzJsu5Q
xpHuh+z6ifBZuncj1oOgyN+stuvHDxzwHI6Y1rsIwkhHFL2RKmXrd1niX9PgwfDX
3k+cBQur4EQcoQJOtCG3sZfVWBjCbM2KVQB+LKx/9NC3M0PfQftpQcDyLBX0p/po
2Qrvw8mPfnzfhE5GAZi7nWyXVcRjQP8lMCDiiEOPfL0pbIIFxwAR/VaQBqkY9pig
xenLexsZekocCcKzeRTtPh+wV5yD/B/4JEPPs191UjVasfPiC6cegnx3sucZsGKB
6t4Lz+zVcIZgDW0ppYft8hoL5t1TIdno8GIMTHZ4cR4cgGakTdQp/Q5/MZMbuTFg
bukm+AdikVwh29ZdF2pOWzbObZcHtAYQrNLDIGuJMiVmR2QHi1lkPS32+od9e+vy
3hAXANW30iE0envLd0/Gr23ZXbJ2kvHPuCdTiNJp9xaZ3aVtGjO100W7uOHsK1CC
GqbxLH98YJecpLCsY4XLTaQNVZZ7OvgTPqSjWkypQQzUi3OhxCX3YgUF5ayfpHYN
GlnCTPufWbTGikjLej5lxBBdVNWL/RgVyvChGrVOFTaoHYXj2OOZk68aH/PROfOo
OmeIi31dVYEKAcJ2l3cDfcRxP5E6sjpGHMaZne6NZPyo4c7wiGd51qmabqVZsiac
ygUrq0tZ63siTo3B25grOAgTLGNqonatv09CSRoUkE2yqFT15304zHZgNE5GZcgE
wHDSbH/vPbEY+UsOqr3XmwVgOghOCvMVc3jDTXU/+cpVTICOzbGCbMryGydKhqK/
VoFs6bYOyLdnCvLrDAsYclJzhDEf8cyeCcVj3yqcpvUSu/nF40bcV/b0vCVTF04W
f+ZppXvHTe2yYazgUevqwrvpyfSHDFgiZC8RJeEMSaFDxrSFeD7VNqjP1fr0EmK8
9bFQ/c4qOewUatP4tdfBmiuQpQrce6WzI3KRFUhSE972FUg+Kx8LO1xV+iBD6JF9
Ome19UKVF+9U4PmHSOgMYc2UCFx9HBS+6RTcKXJi9jUmavLQz6RrplyDFi7y9QEr
Wg3gtnl+jGbZomi3gfUkRuozto9wJHMiJmnjURrhARfE2EUxc9ratWgYfkembcMq
ZYYuBkYMhPdbF0hGyER+1TWabKGgNB96+IYj/7yqCxYls5Tb8Qc3K7CwQfKl36em
+OfW37LRLO2V3vhlT1z4WinRZmH1P/E4fMarYPZwLZaDJwbvY6KwDwi3JgGbiX5x
f2l0DuvvZxDnGJkMLfN1Wnl2HD6tpidyPJJ6WlUbLh2hyG/4+271F0ZwlFDlFqoy
nFnqsCu8ctkY1w6W2gAEajO9QD5PgMqmtEYMDyYBShCr7n+De5q63NzgTdFzOLhP
XF0ikIIeDLECZs0vS7N4Qc93He4xEuAELQ487tKa0B5iS9oQZOjQiEODJAhm0e0h
JiM9tpVy8/RboiNMfdvxF84yup4pFkZS1j4fmdYVkssQZeb+RvUFeqvyhAaAkTez
+7TaaWO10I2W94aPGbyxf8zRQP4F9GmFIlETYzLKtt9W2Sbmdqp/zLTGiTNlrxc+
CtPs8zC3CQ3YNyd6U/iYPV45RywbJVHSsr5xQUrgYVgGxIVrJ1YNEoUbVEbTEb8b
DMBOTAhjrxPFSqqEikF+9tcGzVg0zi7eZSAfdzOGwdlNjMdhl3FySdwwJt4OuQJ9
PtHDQGuX7uPwdLijXxPHNBeJB/Tmcw7SpxNDK1/etx/xjfp19MAIMIM2Atoxzogj
hLSlf3RwlFWkQ0Rd89PZ0X02diVsNtHXdRbhChnOzpT7cnVvkpbKlskUtnn3eDmh
P1qWTq9ic/ifgRklRB2eYwo6vjFIYKj+6zYomVWicnv++AD4DlDGi1w2gLoZYCfR
0L9ru0IO5oLvbz0DlYoSafx3BlVqOJuajO7iNa0TyT3q1rUThY5+yU/dAU/8Sjxu
Ci0jvOZTeQenM5dM2GfnKul2sK9ojdOeU5wGHWIhQKrxeG3yBLm1u7SMqLC5YxAr
pkFtB7DGEfgZTjamrOFvjm9rG9BzkR/0QPgngMvKpu/s/OSWatTM0jEM+xmRvBtO
oHUp+u3Jqf7QzyhXSP1Sixj3HNt1tKViTXCzFFTVmQVfxJyfZ5Qfk7zVBpikEj8o
wKJJhr0bsrR1ts+KGIYtn4Lh4bTk+L9dw6vDGBkPHSUkXQhjcKM2UqZi9QHJZO56
C2wCr4gKqb6dYz4psHy7PVHKZ7mkec5JLdkJBMEE1Ks335ME/pK06I7Q5ZCydZ6t
BySv9p2oTl++fltRcKduOtv5uk4tm28zJdiU0nq2dYycffS34fJlQKmn51p26Kbj
1tCnz+wLoZd6zUHX8ZrIToBFA+lcGGjGcN4v/HDnkipNTsIWSLZU26qn8QdVMFQT
2T0m9+z7TJdL8KL4xLTHJtzDLvKqdKO6MnXVSBSV9a/Gdrj6ne4eaZ/MnnfPol7I
M0/Vka2dZieaYeykIQNIgbq20dfHVSMd5sKevd2JzqOhrCCT+bXK/vD4AI42S0Au
2rx/pJTsUVOUu0Q84mqhmXf+udrt8AxbV2LwuV++b3jsMCwpC4v9lSm7tC+LhtF8
bkZD2F7C6JR/6ggtm7hY56kjcnzOvr3PPNtVe/uHvanWYNIvp4kBFjUUaVMn+k2G
yd9gAFv0JeLwkzXRPhgCybhUaxAYHdRScztilCPm5df4/Ov6WtpDiSlyAGqS/R8h
LBkcJAYV0oHdZcbCfh2EbnrPrObc5en1OmhAYciMLS56wKUSu6bLdIQLjZ8uk2ec
Bg9uaF841rd33dL73lrfQbInlSkHXgP3m537hQ4w7bhCshbUCIPO7KvczFF/DB+p
phuUOwNSZsZLc5xVrJDNHrV+pKM1A3rXkMTcXTDdZP2UxlY2pI+1hk8u2z6ONIuG
bwBm5tR4XtOCbmy72a9lPslTdBrDtE7mFKuL5K25gxx075UVR255kdP4kYJHikxe
76WDqcRbyAYDlhZup4pmqzyw6f2BTiaMmD7hrd2s9IycveYvZgfhZygZjf6h38Iy
wh9bExMVjDaN75m1ZRTBDBuRZYNwjOzEg5ytBxWFELR0JE7tyntjjbEVNu9+qhsG
A3Ej6GMcGWOJxf5DfmRCIYyzf8FqP32wSLo4zfWt6eVYxRFEJTPBIWlT3MRSO/5a
l8jhuvjHEFM9HP7f9kKuURXdAiiaF3ovdkHIFxa4773Ja2vlGxycG/MIQN2F5iGT
+KFrmeUvYkl0lrfwroLKNSGKh+jVwmQxndu5S5CEqHHHWJqTxWqRaJEUVlRHy79K
u8OS2dbJTmNBDBQ1pV64HDzSYvzEppxvPMZ5fSQ6uK7TPAVtrafBaq243kI9MvcH
l0Oiid+w/+RRkwW0/j0kNSYY6YKsM+g4rHCuQ/XDpxiBpiuWyhCn9C2CbTAzopRe
sv6j0hR9gB3vpu2LYY6LCT9icbO+P4xa0688AQMx0/PyMCp2nzFSVmfIcMn+pO4o
4s6zsuH/EzsDXIeoAB0k7T+lm05s3q+am+kcMrk6GB3XxJUahdqdg2PJoZ9JrGA8
ZcaPpGTd9yn/mxgHhdDncmVR2yi2o4GqlgGrggUua94evhr7BPponHvUqNe0GUfM
x4NRMV2MsNKdnkK9udfzfRBi0no3dQ60cKYaegThrmneJc/y72I/ew/ElX45ZWX0
N3hvffH92qWB50XbFsxZSukk/1lEJqo0fFx3aWX4J4bRseKfeutFpzhQCy8bC/y5
NQ1auDlNBF5igSnxG5X8uTEV6eCLwW3yWwKjWwttnqgMrSlXuCfJd2Y2sE8JoJ6Z
sBUg4dZXFRl1826ggr3KBoGsrlFFMnGu4WFPHxaTkjKHSJS3nWB/EW/XUn1x8xR6
ppyT2KZe7HGgJLRsoTnT/x6HOkNgGcyb960gADG7rY0G4WCwUSGEzD+MqzJdPJHM
d+EIef5PFZL33HKuaDC4ncMy0B3whHcyvSS6qFiF86DHwX2N9R6LCBQu+jg57kWN
bImlocgEai8lDsWADjy+iugnsvaZ2EFR7aTCbXF5aVyhbllqZnoMNFv811bU0aRp
EqIce3jf0wKC+SsoMA+eZ3dj4AKspVIrvADOPryUQhsTF36WvfyXhvn+g7oxqszL
HO0bZyeowGAgtx74xAS0FNzRqW9w6LMdmtQV/8CJvEAXfrkZSMJ+p0kZ5/6q8GKG
XnH1UZQoAImZ0lbym8gRYltLK4FXqRNtAy7G97j65k+JLffXSurgDcXqfTEnlx2G
ikQ8PkIODLWaMefX6ylMwXb6VMVP1dKiQwtqjWqb3kvfs9aOJPVfFDVxLZgzuSC7
DDDrrMJJuBYEPqBASAcEzFYQ/Oe+7qw4zhNzcmgXY01jNfFA5J3YVhIiEd8R55E2
9SNfHd1Yy5RGVnC9s+PZHVIbFp77tLPEv1bbJnN56hJwFLniwjNJ7/QjU8RFc1tD
JsjFnNJrDlNK6BUJvEdTdZ3GWkdDMRv5b4rknqYiBm2xOc+Ill11GpMj0AmZeLk4
+xFe0QDLinjVfv0b8uaIW/gUuQA+za4lFAXiuMW+3IAgSWFcsoqdEg/dvg8GXm93
dYHOW1ktk6xiX2cPmQaRaZlpUYpWdkQYffiWseA+2zSyXg4lGAwjraKAkyZ8X3I4
R3jWCVPmKq08e+S9VPIG0p0mKf6NrdBJUDwXSfy61Ryt5aW9kolapgNPYqt4soV4
0kws72/u6VV4Ad06i1+07Qj1loTyZk0/GCzuxOJU1ZUFX9cnFSPUQQfA8y5U7Bm4
8o9qBUDVC0nRS+SaYtlfdc7dzKx/FYaJ28utnPH/sXk/EtXMRYRHbrvouoAassWd
WQAtrMpOTXIyL7dzFsu3djDQD8q/Zm580BakmsBKK//S6/G6fjtOuPuVZThybGUG
9rYmgTDigCj/4ast/A9ynYbno3XeIIK+EJt9igNLrYsQIS0agLmLh9joIjRoxmEw
MckRco7NwyNPi9CFPye9vtDt+J5XH2lkPIzLWWBSH1ghlBfiw1OHz/CsAZgAKKmx
vTa/fSPpQccrGef6EVJRw378OJDuIHhulfJbWYT37N4LuZHfZxuZYiorUPiSpX6r
MA8UYyEwmJEKBkOnjransLsKxSYNNl3JSk8kqo58QZ7djB8mwZebEwSLZehOIb/D
9rIfE2yT5chBlvSQ9MnFNFEB7ld00dpMT3LkhymwYY4KiyOFbIJJ+8zRpZ2xZ8aR
YyVeUs/ZN58zxojMZq7VEn8UBioqWfd1XkA6nBUMn4dTlU2xxd5LDisG2nHg37QB
MU9/7GaZOicAQuLroMbxPLyh1VCWspn8OXbIBcB2Lyt5LeEk6/A7HPxNB9/IMF9F
HPFbVDDc3h7oRwHta/NkY8lA8wWQfFr+9OaV2bbrP8bc8A+4lb2mnQFRWGo9EubL
Qc9E9kQC4wfg4V5dHOk0y9dOhiorcM6xVPh1qCa5tGqUIoxcjOTFQ0IU/z1AMnZL
nFr4hb+NLNLK/V508sYeIL0gCCN9RD9ow4eoknlXeyK+zWqzPCozFKN9ECBmIFpK
XZ07E42UZ5XPdG3yN+pPhaVvSGmuSf6eRR6j1KodReGPvWJ5Vyj6npCN70Kgme5i
qlwR0h+y/SEIEZh2AYTyep5hitk6JLYK033yKsRvLsA1vjw+KqTrV0jmWD0GIrPJ
1/Eit82LIyke5gSnW0rGfZ7Mey6gAVAVabf44xMdWEHTSLUtJ3iqJUC35GEvr1VJ
n+hHMm3u52OVYS/mPw9ustkvOsDbjrnIKshXZAyk115RAhSgCU0pN3yeEKXb93ap
oFOlbseUKTkYRnjFouTNVj5bLOutrT5HwyvnzzNGSJfzfMVLGkZrsPMrgbwIA+0s
RPdFZR+/9uN4OvtJ22nDq5uSzhygvIXRIc357lS4UOlb7LSirtDiGkZ+ZvcYs9Aq
aEis2lFmxFxmJUbHTGk2W8KACrhnUxo6Boay/BvVLtPFFI8unjGQEH60u73it5ER
d8SKjPyZbKS2Tl7zNhEzidwosbjwgzYChTjgsOal16Nkr7L2gSlZuprAlqCx9lC0
YOWrHjyfy43SgAt4nwZmYrIhSt2cgmWKcTvEudo9MD34/PK52zZz7i7Q9UiYcWiz
J98r79aEkMZHlT0Z4vvuLK1aWmYnntLvTKcCAeZONmO6sJXZN4Shwefj+K7M03TN
EVts8q3CS+EFxyE0Uq7zL3wBHjQ0o9xNJU2mmwljP3yU9dL2ObAXDgMCC/1c82R/
w1TaMZj0xRgEai2XOF9aoi5OEm62QGVNAn9kvVebaFu0mane7tiyw5kDAYffdgKK
TzKrO6/0Wa4aQbMcamwIXx6cUq72rC22Q53IZfwaocHEN8v+FVtfBJqHlh4dDkZ+
Yv261tl42zdi24IAG2M5zLcyugAbX3GOpYKGl6d27iVbyPQEUp0gTivHirrCoO/5
dK26A2zYL8QM+z8TbIYEsPUQBF6xmyCZUroVQ6dMTVOjG2TRcOLgc8nl5BFxzZtf
bTAFLQy+i4lsDDqV5W6VN9q8EDZV/TlqZnBRCEgLe2h5j5XrLwJKtnTDXxbSzTlE
0APv6xBHyYXsBb43DAqdJ8Ac3Y5W/czpwyJXmBQzCd1hhXA80BV5dr2KyKygY/8Z
5I5KHFDd85cIh1Zzd7xHHV/L0R0gIIgBxiq4hK2oWsWkj1A/BCl/CFMlrwaikC3f
e9a8bc7EhJHWqSZJI/XmY29/s2fGfTVbpD5Hnch1dj8q/QXCF9EA2bY94ztL9QMJ
oc7WmNQE6oHYCPo8jjh83R37R+dgm9dVYnuxp8EyqVxZt6Puw9cR54QHZFQgO98n
blQeszHfMTnwrWyGYfg97+gft3S6jcjoCcGo1MdQeStNYeunQiYJwDl7zthrnVm1
H7nR3UAUT7qbeIKOOOl8fWG8nU2GM766/Gpqv2tku59l+un9xQxTLANFsmQRELuH
zN2T0cHujtY1EZkEp4MNRt22FgeujvOGQmStmy7dSe4qGvOw+xTRJx2pqjb7iTkd
ABoQUjEmH2HN0JXxayl0ZwIOEmTqv0aqjDywxqCt2FU3hvAMNmyRYvJfzC7nhwFK
gHmTRl6fi8G4OpCybw7xCt2GKIt/29suHnDY9iVAgSvZnck9a4U+NbMY07xFyG1h
FbklOZzT6Tb1BIc8JYCLX5zrG2vYE/woickrHP2RK1mNwSTOVJg7ZacvKguosXzs
je31XV8Be6UABOAvDMUPxuvc/Cce9n9D0dz3qOxJKHGQyTB+3QXIE4LREG43Cow+
2oehIGkXiEZinVRjyGN3zWGRsKPRqZDG70cw2nFrvKwuKsVWMKp3yjl5RWMR1itH
vVo0QZ9oXnBAJaCjjPqOwsT8IsX4Mw/p7Vtq0wZ0Ziq/6cB6YJXBwuNpqcdtOTEW
He1ogRVuAdabLr11tR+6oxgXZQ+uFNu8Jf8AbN3RDEziW1r+aoXYa5tq1FlPVWyY
3+mkmrZj90XHl1spaYPlOfQurnsRpilNhpHvZ7wQSSDlC4eay7JrzTfiqIhjUznd
i8EaIb4PeF9NsBPs2WvbnEMRX2gHCrBnq+BDoM39Egueefs+PhzEx6juI+MF6fX1
Nw6FZipB1O4yqg1P0H3/RFBadzl4pE7OBMgNEW+h7Fbkwww1YQ+IXKlGSq5FJ0wO
7VDj4QjmvlyS3o1hR5hhrxylbnW42MIs0PF7jlXn2St9DycdOltnr3/BZfQLHiOy
cThjgBM+WBswcCe4ZRNGsEjhiLWHtu7gwuet0Uk5JEa4u6xfNh4sv0skLqS/GKTH
hdGzZxo1WrlqH6Aw10RIs+yX2poOoKwqfV4WUcU4Binmgb6JdFQkWtwlBJWNbLJy
XWBBjMPrD91Q35cmJF2vn0MoWbpZ39ohqr5tErdeu2xJsaVmQp0dwx+S44paAzav
aB1rTAWZ/YLF+3d3BPT5DDLPcCh4iW2fXcsb4v4+BhbylWEnw/vqG/iy3BoVaSeM
h7yG2f/tKgqjtzGUxTdH1klSsYbdLwIeMOGeKn4/60dt5RsFiWFLQaudSCTTVnWG
Qs0WcW1hCvVcBlGQHgfB1nTQLTisFF1rmWQdUpieMm4W4KWid2c6XgQNIj5UqKzo
k/P1Almmtqok+72pqmHSTwUqP3YqozaAtgj1OBCS1jlPlNsnB+zt77jQaWPx1XME
jLlguvhonn+JnZ12LpKzwplSrXhnaG40FgNE4n4NwLmVNgECLiL7yLmH2LW8BGhi
DC1PzeA1o+gt4QNqXiVJXJMIlX+sA5eZ7sHB4QLs9qdi92sr07XbyQHDZYvfCCnz
7fadlG2lXQoURPEtuFOCfzJRVjFfbSxaWXC726datYym1TbrMEFm79FbDU6dNTBK
GoEhpOcyPM64q/AU6zYn6xQ2xoTAzBeR0vBtvH/OvAArlgeazIawGIgfpQVhdc3e
O91r7MH40y9V5pyh1rDDxfYjl3xbZNs1aAb2Fh20g3Jkb3MW1DFwmcfNmZf+1ZAE
eaNrVqfleDiH3I8t2JUA+oe9KrZ9XDLdG02rDruNAipedl4q8WDHGrDgkTvhtwx2
KLbmhjj47iFXSWIfgOlif1XnUzx5RnTSUk3wTNrEl8zlUXULxTiG58ik9T/6NCKV
jJQtF/iZbkO6SLPAu8L/KSUYvmwRqVOI9W98UWShyFGhbuDSpgBK0oOnE2bQQDE6
+GCKFVldeof1aincCKXz8qv87ssSjjrXIEdtHNo3CEafW3AknX1PL2+NOHuiy2Rt
+FZDCa8AZACGJlskjji012azpVJmuOloxh216uaK6vAwB+z821CH2Z/7LnfoWBKD
5U2bwbPydNoQGB/JO+vq0/qufiXPt2oAZt5mFLmLuk7FSCg8g8vdhn+Q1FLpVHG+
olYVdBT7aso18Em8LvIqBWxdP3V55WkrVhxBPv+mLsLTAWBIMSrv5SRYxJoUOTkq
cOpiOohDe4vE3jaR704N9+umejsxEYAYCr4ykfUOWuQdyYIxwW2tsfXcGaLuWFin
9B2Qx1f+4vGYy+0u3Ni70GvzSFZ+QhuaiGQfywT61FEQsCST/Y12HBMh/+nb+wVn
gRoAlZ4CJGkMUFHZ43EUM4gZt08meo5Kd4o24N4GLKSwClxKEJMET3giEX29AVqd
pPKsrGmx0Q5HcjUzuIzIKrU5f3EF7LEYqW4IHTEoIMRV1/PNYyqX0U0CVZP19Bri
QL2EVvfb+/hyNjbhmJ3/rLWDxC0uzfddVMngsUog8b14O6fBEK63OAEhxjy3Z/C6
o5ZrJx8cn+WmFlknZEm+EseSqIqCNF5NPcTVHiulBRqGDrqLqsI9+o1pLy3mEvzo
IQWBsa5ZYtGv6+/1qWITz3G8j0toCHz4J0OPSaenaWKpqT0K8Pt1XubgELUe+KVt
xkSOWTXvgN/eNBbV7xdAiO8v/x8ht93lh/TDgTttSzhAG5JAJEj/JTYkaOmZrJ8x
LYRNlEnSDW5lksY+9tbe5WQ9SWM9PRhxOWAYgX26CVVmXYVoSsC0MpoNW233nhbM
8uIcLSLgA8/zjU3iGboEp1NKqh+/32UvvURkW6BII1rHiV1iUX82sXm8zjkYDl65
O4f5gBynr36xHBXVBHBvgZ8ckkHofPQjfKSHWdW7fGc7gLcZPsSSc0mg59q/7XX2
4Zr0tdjHzV5pCQrkhLYG7QlXJpmeHFQjc/EZeRN7L340t4rzLOYmOrve6uKY/EGP
mNTXfPQRYt5Lprd6NuPyDwwlmR6Vv8CN/ZT4Ya8TVe2YhkjZ/YSuH9f6i8xEv1s7
Fg68muz/cHDJGBmZsUcc5hNXpfJqCicdTagMM7+1/TBpLBI9FG7eMRapujoJfZwm
4z1EGN/etJ4tf0VSEjbjeQ7Ek8TdxrguJ0WcLZdVGRaTwHEEtrTMrV+rAscjnQ+L
4me5OyWZZvFz+sve7DLpDMp9XOMhQycGzpTkl7fuTzwdoH8wJcMAqPFU92/7kQ3h
s3vTL3RBR1HFljFlAiTBcmz24umO2yHmEqmKlGmnTzn8DkTUGZ3NWUc0w9waF+sA
D+picF0O1krLOEkHgjKxUsLB2I2FEkFPK2AJkePn22OWkiujdOfSKkYMEcm1FjR2
kbVAlADF1IeQE2dK6hyt+eEbsgOhDrklxX4SYKpXpco8kTo2ao59xPOaMOpG+koG
ZUXKDgriICdgYkwp1OypAEIfHrMCuN1ugG/QbXyXFtYoIHQwMDDHw0mpMfXv3iHa
he/4l/BnHecGqgV1y149biozih6w62DoPhb0J/aSmlH9cQi7oCVl9LkkFaz8Oo/1
0Utm9ZcHEWem1dnEF3DEYo9G2f3qd2oEaxJKK9XATpWAhv+Tyl6dmm0QAN6olFiu
uZvYIRJoO0BlYgXN/fzMRKgl8MwOthSTsJ4lZa6d277NYQJQdc8RF9MPfULaLt5g
EuwOgN1Adz31NnKUKfwVMZpjq0QOYigL+nOOzWq6MwMZtk6L3CYxCnCwz28inJBi
0NIIy4vEhf6ZsLVO5GBPsXj2FSeea+HrnstgnFfGos0ewn/lpfRPJpqureO6X7CN
7JzZDTXkeDPbiSROvNfgkmmR7x6i9z8cDHYZNj/BVlbC692xZovC/GevrMpvUUzs
oZYMT7OfymS/lAgWKTewHs2ukurM8s2E0JynLYYVdmox7aFDTLX2ecddpKMw/ZDc
mpDw1fWiUn4BotVOplEoRF4frYfsnV7c/rREEWgejfZODbbdYWZneAgumuUdH4Vj
yeqWoqxOgQ/FCYrGDzW5mH8Qkzvk7tTCuXjC/Q6po+pRpGIgZL0KwunmbLmutZUY
7WEFUZ/Mc+p5DrI7ameXETIoVw0aGTnJHCE+2SkD6kMu9tg/LrfSXXeUy1GvFdEo
/l+24fM8QtXp3UVOZ78cB0NGMkQAlSixFnD7ktIvZNxoHgSuoE2ERnM/ktFIetob
p24vRlqKxL7ztgqHs50b71lZTlN4o6s8BbxnGgWn++jWNv4YSfklhQinedY8hAHG
AT8EKaqYuprCIXaJnU36sHZDoVSbdl4xyu69o+EanRfLPMWaPf+oF3B85AR5wqmm
Bv8Dc2euMF92e52YWO+c0kgxiP6A4Dzq1b0ftWupIF61B6UK5bvhn0GabBDdfxOh
bhlk0cvU9vHm5MKT4ryVuXIXZtS1wTisZhyx9EIV3GysZ7d3zysJ3Z+qaY92VHhn
8Ibd0wyEk0mrMIqe+HvK7zZuaFN8b//VDKHugYVYevRFWIMrXCqOO4YFsQSl3dzX
/WGv0ra9Xg13UVfniQfFLpwZC/ERo5nIrSR0OY+89z/XUXT6zbLnWl8JGr6dr1PY
tHbZPC2XCPK1LIyzWLveP/ZrhxRNNgyFRzjdS5Klr56tAuer6U3ba2trCGJjsC32
r4qv5OQUZwTH3TLrbeSXi5fylyXNXan+DhJ/BU5dRkbagnseZN0K30XIDH9Qyqh3
szRC1C4jD9ozQGwge6E/tBG+as/lNFMygqPPRGMGU8MKScrIr4gHbONKEzFQolyo
4WASmeMS3NaJ6Oy1Is0l4fqeHNBV2Cc5zjCXwMcvthOuEYqt1ceP/4k4Y+GddQKZ
uXowYfAD9m1uhflfWLo3bQldQnDxcsSyEBGvn7duoybdiQY8GhnbWSwEBIGzRrH0
i6W+1eWxJ6RyPeupHup1y2acwvwRmJ/g/Imky5BKb+qHUFmcuUIDiV4DXhgmfSl3
mXqIW3B4q6TKhJzJFEFD9h0ZkJaYzMi4AfVL/IRgcZ3Kl3BrUjchuTU0uZ2xXcYi
pNTVDa2GKoqDpfBUE7jukfDJ14JyH0/gAIHJv6AMb/MDjnw96dzwpEkhPq5jaCa8
2FYE3yrgeK0WYqrBvqZ1HQWBzFLUpy9etFEzaInLo8rYMIBx8Kdh9b1y9vCOAR42
imXfAlbElNDGrA4pVPbHMNAesT7CYic2YDxP1MotIG9rFxLFpdJcDtmyny3YfOIV
YwJkku9WD51YlDnFut9b2hNIS7QH4C4rIlA5AtvRZpvVpmhSutyOvTklhNMxgOFH
FFzVTsuBrQBEvZJ4lM/Y59HOqwa2a4HbCTc4Dv8LGlyYriv/kCA4fzUTOpkSDMac
qxr4GI1nTpmFTB5lylFPqoORzm+7M68CvDj0IrihFReCvqxAva5C5LtptFHwHADd
npIMkD5JSv+vSGZ1FZa6TycMuazWOZNdS/pdrdjAMUlJOurGLn55+KtiNkhaEBJ7
GTd1wyoqyZNt2EayaERGewXbqMIJvSWzSs642TD65D5ZOyWWwgFRJSqqNxHi9L3I
TqdDiJzgWLV74PE61BRX2auL/3MZcQ4juQgoo8R0OVbd0a4rlZMgF9pkINjy4RBN
0Lq7wysa6eHPvxxpdaLcbLE7GCUsmLX4Ip498C5JYY66fFSv6GPeqU3Oq28fph9V
jGrUFfncRsuJB0K8OR7uHa2jF6JLBNQFgO/n4+5fm4M0fyGXDXlO1PUe+cJxmakF
U82Ji8SZFWrUfaBLdzzOq6Ly/CfAbUafVbEeAxna1miVSrLr4c3lmTgau3e7LeXa
q0TicJ0oTNe3CxcCxIFkiXrzwzQdir0vxXjkeki6qUfWe7Z7LmAPDnvwvvg0cB2e
skjGTfgn2tT9qcgmSRt1YY4Kvtfo/EfGRyZLDmGunN8m4WtItYp3tCETiYd9OiYY
8/tKx0jSA+egXzYi7JnhLShGKZClM2UCNAxLjBTJjLO3yrH6bO5Fs3Elzzd/9ZMq
VpaLFBUkeLMQkwrKai8vELwySk1XgkHMDV/gwLvopHA6ei0L7SH1DyJYILrLHY5J
KTZNytPd+evpo8n5XJQgT2uE+I58vKqwTLlkboOZvpfP9/dWBMP4T+9jHPvA0PH8
ojOIayCt1fcb/jARaZmyQPHU88Cy6nJOfgkcIre8Btt4lqFvAf0dAVrOIrSSiDfJ
7hVLl5n6A7Izp9cLz5lW4eDEYuVzaaK1XprO7sd+VGALABR03UiiVboUH/o9f8MS
F3HrzzJCXk2N8LlGcIzYMz9qIykhWQrPPPvnCJnC/Y5wYStCN0P0MVSzo0kJhSGI
cfUBthU2RcIika99jbg7LkbePHKrQcLX1sXar+xne3vht3BTkYHYjW+6QyBs6pRM
GXPTx7T3Dvxk9JYQuoKNet5xoaEVhi1Uu+AUkY6HY5NFsey6O9+3qyFqzZwcSd1I
ikGBrXzaXgcTMLE0wCan7jvA41tfz3I7wjrwyEzVqe29dquKIy+BEN9ZPPlT0k4j
REwnmt7QbzT7RtMLM/MBQzJ99m2uawv4/QLgm88oUhUI5Pd49sN+v0eeh+vX9CZ6
dDouhEY6jxHhvHV/e4ViI3FI1Iij9UHa2l5lzupGQ9tMeELxZUymqSCpointqA+z
IH8P18RmyY1B94RYA4++rBhgbJN3y0mxKPqhv7Y1On0kkqUSIagSW5XtVl4CCwWn
2066InTwrq6LUzqHnkczfvwRRtCjP+gkmRaloNaB1OOcOXJLmj3iC9TN7T698D/Z
X2d2hH7zzPEzjxTOjcWa7gFjr2ee5VW27ilV1LeTs9cBITTQ6ekZmDV0F7zlWKA0
83/h25aVQA/I+VAPBucZh+zHPnlvokJqQD+6jW4lMOGOI8hNhXDMHsgytVXk/FK5
zrgSaK/mznsBv2HBIaUyFg4m5rce/m8IxkV8H8diSYjL02cFwvBntQ0v0cq4QKG6
IG2+3JCOK/nnaTFOziqshnedcDVNyJdEspTwMMDuLp5LqWIGT+sHrKidNwJG1oMd
dwSpjc0iG6TzXkhOckYJlfDeMXqTRyMq8/gQiNCbyrHWPHc/6ICPCzmFxZDfgLFC
yhKosB2XQqqk1MFqyNW8Y1JXZrJVGL8hcVA4G58+eehHuELaA3bDi07ez/GpTto+
hhvfwN3Nlk+2ehcFkLW6rnn36V1qrzp8lOw+dFPVZ/CjgtOww2CH70Z6aSSO0x5b
D/1lu/62Wv4LSsths/tUtXoxZwxDgOmjpL7lwSSt9v8Q8E+yrgfEF3R/s87O0UDj
7IDUse1liKBj5XqsSdQ+je9IhApCBnzI1TDV49hkQa8eec4xSbJ1f+bRdNn1Fq65
Df0ZieSsgrmaKdkVioPpkMwox73uwfVg6C+2CVsveoUBAeaNlZPdy3dSUiqIVVgS
epJqMOzJWC0cbjqEeedL/aeIRHFdM3QQyydGfRnA5rZVjboOcmKccfEg0icYyICP
jZ5WfWutqROX85yh/uD6Qk0QuaUOVFkTtmDIUsD9xAh/L5MWqcj+ArV/XBqSXMHL
sQgqSznOVgJ0cirI+whL+ychDOt0JefGhv7OJ6m+R3r/76NyB5NSpbqaQ6NZ9LOF
EGvSnVA+vIumvQ7ua3YwE01lzmj0uwyi9SY7yoUM69+7pJc1zuFSVe6HfNKxRyJU
zRaUTXCiQ1+RTX/ZpIljjLTtRpYsa8BZNeMOESpQG4HbGvP2ovqs85ozSavDNYla
WBA5y4o3rfKWjy4NKNZq6YOcs7bmqPd3+w1XGHyK3CZvDJVUGJo0fVTtxbk36w4s
GADLeQJjYQiHZ4y6TJCt7AUIIJArEo7JW3zNEQAfX0Sbnx6CwCHKcr10lD6CQlD8
ThixgFL6ghzZi2UHgkvtyNchhmDrkYTD5Q1Qm52oiaPSaSH8vvfXAnWZeNEmLw3W
KkAvuPQ57hngTQpHumfdHbNZmG0n6dxFYWtCmidwA/uAaRVBJJp4wLjPNCKKIus4
vD7RGz0WbjRco1lyHEwhMXI1mnWW7Vlr3tet06EsHL3cN2PKbofchcZh5h/eIbUz
wOsSS9Bn3iHI+oLqxYoAD8T6MjHMdue82ikhmPv9ZRgAqdRWE2UspCHcyre5Q9tz
EG0W0Ml51U1uhGKRZ5OhK9RawsH/wRRKpCTYonhNxIWkXWL0UkXae2smdPyfDRBF
NhEJDjqznFkABQWvFFrkLHTQKxZ2F41nb4N+uPkFH12zayESTioCiXU7pMdlLSxi
MzjdbFqGMYFV/7VES8ylELO3NXEUNEgd8sRanWyLy0JaPe8Ecx/hCypc2aeTD5L8
dq8eq2/iyuIQdKy2qQpquB5gltyp3kBGYkhRYlgkfWWWxa/zTIi/uumkggCyGJTk
w94E2bowU8tWXEJp0iViL4KdJmLJaPwK3AHRqECe6fYiOKCjCAGgh8e96gqO+Bng
FhnDyR7xLT6Yoe6L3qJaaC+i4GLsR9VTUm+HBRJ7zahf47aYbIE/VbvqIj423O1g
CUkRr+wayUvfYBnMlYMtWIa3DKKhvBmz0oT05tAByDzed0ydojjD0Xw5P5MSAYMQ
n9cmpVerJVgYn0RIihlYTYIIVogPGWyMStxbABD2acXCoIFl7vkqsB0ISFZJkYWg
HulEC+mygrXHcQDvEw1m6dVM0TvrVkyvtHCh+aXX8vJEUPEZUmd8KHWt09ESjUez
szC4T0qz6VmwuF4lc972FF/S9zY619RndMUIcqu5ArrMGFZv8DRHYZXc1I61dXNS
kNCLZiBP3EItiIEILp17I3wIkZ4YqWljD3nCOaQgFrNKw6hqxa+0ojeDu+E0x2JX
isN8gCBBmPIyFz9IpSLBtICfBFun4F14DqwiXiX1V24i66bI2wRfjX67yCMybPWg
KQWIpToBe2NHL76LYuLI3WQLkHrsYahvfhv7B7UL6WXVClB79yw4gy//CbQn6l+S
t6XwHvzb65NAUGQb/kD6qHYtk3bGET0rAZ+yUojm96xigD9i0usUo/gDicwAIzGa
me2mWx47LRfeHqi0lwbfaulLCoexUiOfrKIcdJafASWImAEAHvmifU2aw6TV1Kql
puceqjzv/LvEs/yRox7qSQuhLS1VM3h8suBFTm/XnJDTA+w22Gdq57dH5TK2PXl3
j0GEXb4nEq0YuEzJZSMqhFwjKhRHMcH7XLwH2wGdgeTeZAJ+dSXgNpLvgqY9+Rqq
oLy17WqjAHusO2C5m46Lsr0JMr4cg/HG1/j1xJn5iEVdzaj+Y4hgiyZUIBOniAYG
GKi9/dfJX3HZ8TXRtJL1aBt5puziAXhPbY5sSD2l40YzuyEBn9wzAxq3mE3vdjsR
3hsYw1WygN5ebTlC+yGgoU8Hz336xqg67q/u16uQYyiK7mDA74UqyEqdub/p1Bu2
O0yk6ludssaKyADlZ4W+wc6+eofj3q0P/6XeAbp2M0kIVt88U0GgW/wEbI1Jwg1y
LiiXlY1qxRSnE1+uVdxqNiz/Pjy/mcQKADrwvUGlbE0PKR27tfUgQBrp248YNx1Y
SJwoV7MhaPCgQHt8vAljnvu+B04RD/wmUXmKNFLIYaePg0vZwcCB30qY1Bq5P8Fu
Vwz5JkVKo4fVLse7shDzpJZSCGQARtlTgXRr/b93H44f8rrJQ5sc/huSQ1VRbfTm
+Qm24xkf1g6DAg1sTQqRmo5LCImARxJ+DfFkSGX0Znk7/h6TL2r69s6OQZtFvqV4
A/2KKayMeD6jZZztuH6EuB7U/NQZRZYA67q1ODvJ2dGKgntZYkqg5AKcV/Um5uQc
ZpPCgatBLevc1k6c5fLHBkXSsr40nDEQnJaSbc9+CDu15PX+PWgrtsfn005am+ck
P+sbYlD8pb7JqtXyIHLwYvkCsPFlnQQik14NMMIElzV1+QtP8MEMiwWCUCiC2+DP
ZOJ/gVXjhe8Rg9YUdUFrlS3osGlQen6RGJbxnuWY1dMt2UClY1/Hy6fovu/E+ROR
5vhmijrDhMNW1erNCSCQJXhgjfmKNyUEhKcWCgMPCq9AKUDcC9SWnzr41mM1WzAA
odXHsCyhFZKsYhhimGb2gb/I4MhfYXtxVezFjz6/rLRrw/MkMu0N++PvG4/tvyWI
Owmo0aCqXDnVQ7In9qGWMrNM/KskpFo8QjyCnvBSQo1cymErtFhdiCgVvfdsxvKn
OV8+FjSUyGSklOQjTXRIglkynQzM6XKG91nwAQjS6O2J6U9vimfx9Kq+mPNMgHVr
qpzs/ywRT8zYvq2DdufHZ+BDnZB3aWEcSAeEIY2gyH8I60xiGy8QE/FF2pwHCQ/R
boPHLtok2So3s49v4mvaXowWTtSDSo5YnO2CTT+X0XvWnrs2gTTop+zEPH9ayb66
dkIpsnJrvaqVdGDN48lr2usAywZ3ifvNgNzAo9jF7iutjEKrMOnNsEpaEr2C/lS/
eLf8dRStIscmPr3gbaF0TlPvZsVA6WujeejeqssMIT3ZPgPD3iQcwtfLWBdQZlqe
N9E8vySkcOCpTDToOxVu+/LhIQ/6dWwqQRF9xta03nAQiuOrAwSyL99zSWOnA6Wi
ASeDTOmQc/UxVWLyVrv+aw0AYdrUrF/7JxXk04FNy2kUHH3Dwsh+fyCUcN4TCiN8
iP2D97QTBROtHwFZwovGSDbSoNhk/IWoeYo2mQwmjxHiO9z9IX0mR0FXasT8a2im
vkbkNBqRpOM6XGuz3XW5kSSj2MBeXncMjVVM0jiG+HDau6Z1kHBDMAeZ9DHKgAaS
O2aav72qvSxsz9mCiuoUEBww5FdTgYWZ5UoF8L4I8Av1f6AloUeriqxR3CTzFx8I
WYHXd4XgSUQ4DEWPXR4lrpnRgpnGiFnYN8+LjUe8c35AoBEOjcttDq7dV1o5r9SK
GFptymH0Rn6nPoNBhIn0QaDhdoKBJie0PDkAQojvkFyrSvU1jQXwv9tkCkA1ir+E
FDV7atNDHgXrDw4hTGbFeeOxfn9sj16LelpJdjt4BoOc32Mv1VAik39hrXJlc4kk
dLQAfdTxaeSEujNylpEFU+CSCgnvoCOFvZmOH/hsd4khbZ5SU9l0umZlyszlDmqR
wFO98hML+tsrdFZFFygtTkTOH9awFTbyQISEbBq2HIP/sjK6AmtWR79XbfUgqm8X
NYSE6XK+JRiTcCWyrkTKOI6AiTgSvCGxGQN6TDH71qUJ1f3FL0xaQra5jwiUernB
Q16nTAXGzKCvpz8doF8Zu2zI44ON2BDJvw5OA0TJRW2a1p+aXz0SiHEG7YLIl41n
YwvQ2NmS4eigisyVck8eQqoASW9Ltf4XAPcl7Lfc1uxi5Y3UhfNa2ZVvLbC5m1aH
4dE3oPS1Hvv+afjoowDgBQy3FqfsHF6ht1ERXWcmovCbjbAojEG1qFEHwcDcNyxF
/baTn9XThg57ydkKtErh/iIsAiwM6TiMAZunuUPd61cvili/G3hTw+oJdLLq28rB
v5BfxBeCmwMpRiXl6k/dXdjQkFuZkd8dSGUhe8JdnbxhRLnBNSMjsgMHQFiLf22U
rYTWN+nCgwQwmZDkm/RfeUKilBJAtNjFGqVJ2nyzDHTrJ5LiySJd4GjoySbjrpIV
Wy5U7Pnrmy2pnmWZV1rjea5a5ek7rJFF4fEiM7rZoRbhxRpykVv5O8MA6ia1Pv7B
FQlA3uJpb5jeADFQAU1fJ6ahw2s2prVpJA3fX+GGWbrs1XKp+k92vc6maVx5nz8v
TE/dUZuiqxRa+HZFC3yXsLK0JSxMtvMINgqqRAOctJqRlTb5z/ET571SV97JqetW
3vjwSlAPiUKzMSKaI7kCc5vkeyMyZB4bjO2Hy4ewafzkiHY4Fz+VOU/RQTo3k7EG
M4YPMQ/ejrAYXdgbhOYF37qHQJUK9yVjL+ZfsKbUuwLvgoxNucnnxfWfsqZWqPRp
4MTUsFYG2HxsScCYqW/1iBla5LUHb29oUhWpGSf401wWuEAzRpcAyk5jAGJ5V12u
8UCWaVwguDyzB2uYEtVdYD/OCe8zNUm0FIs2VbA6/v4iCMswDcgSyKWYI8Nz+vUM
5j4P73qOUCoZXe/m8tl7Uubx89pwwL9df/U9pYeqY+jI74Hpx8y1mCQJUnUtw6Lu
HbfXzpwSA/1DRHba5Dv+OYFwpM0l2wt797tA91bJchR8hTM2HsNW6uKzXDQcJKst
fasUjXF1JPXV88D10OOApy5IkpRA505WIyZkB7fgqURphBmIzYYH4Sdus2go1AAW
Wi8ClnJdBT1AvNsNKUKG5/S4/9K4vKPr4WbmCHhsG/QdECK/eJO/hrb4ATv43PF+
USL6T1vjLiWa9Y9UywIgKC8eT7K+ZtFlib55+m1MOox/jTnSx9LAHHwkuw8Tab48
oatCMDEkH0NPfVrXl258QhTkw/SZ7/YzzagCY/wPBIzZzd5so8V855LRszE8RAYI
AEokRopCuKiTldKVjKinnLOhbHk8VYcqt0AA7EuFhBaUZclpB5sMYreqX8HNdf0z
9zeMNBOOB4wWIqf2KIRFQcOZ8WGXqff5Yxifq+qUeNQhyiJiEEpNQuRK7W5Bcs8X
Nflrzvlqa7rL6ea0cUYIHUEGI7EuPf/LriqptMlIAtPcroLrvcAVwGuiuDwKwnRI
O63ommrS5m1hQk293PvNH8TiDBXYVvW9JI/7hGeszO+S0LJ/zcSY2gi5yNTrTrff
9p73TkqeYpGl2zwyZ0OUK4pUP02mmeRviiqy9heiZZFHvms7xdF2p7z8/cYX0Dk0
VKB4+WGD5i0kNK68CTANgt9lT13RRqOKfeGgoc6uSzkDo6X1SRmjl/Vqdqw3fZxh
81xoXWo3nN/4nSrRlA4IOr9ceyeABcccH98JRNgj7JYcpL23PrBuJxJcZU3o9n6g
2Wp/bA0EQzTCipPn3fsToF8tI5WuF4gR8kMXAut4CE9DWeWWfTWc+/mCbcDqBDEI
hs4V6W4Julhpt/kJdqJHsEXRIhB6sMbTjnzYDPOQphPXGFPwBuPoVCUHcocNFQvN
zD3W28TZXYarlDXfy9efNIUebeQrlSMYhjzNp4EXIKBgwAIi09QM+ALwCSP7DTTs
9vFyLqbYVNuX4tezVXBPrNgV0zHUYqyCFEMm5TTV4HiqTnJ5svJwK0pRulA07SxG
DGxZ4HehENzeeSlEC9i1aV00z4liRp5Y1DD2DdxWeNwqCQJD4pcjSigqKyzzzV4N
1MMDwBsV1mex/wRp2EGRdNieJLhfPuDDuu+5NmcdiZHbxzsZYi0j2uBUxRx09VE6
GC7Kxun7/kSRQsujCrBqaDAIpPjJtsIrXf4o1xzuky4DzC9qFbtVBXDNgOfMmSk6
6aDEj/sj21aiWT7MpUxxMNPWMj6Ljmv9UyFlpNE0opBL+F5zuQ0DNptxsC5SLA9j
h6RRtXpFhFLgx3vfx5pTWd0TSUN/CH/fa2EnWOl61obDE8hCu/dWys1KKrnBCAsl
HUCe2rl5TcupAQEazybEZH63MdNQQoBiLh7MdQokvCqAVD9P4ucyqffbcz1KyhLP
MJW6AdWJzXnn/3Addfs/ah0EUZMim21F9vbBp9Pk1HImxcxVcQoPzQQNq2C+JPUm
KjKOh0VvjIvpIS/jdt8jyMzjHzhDukprHsMe7EZWIQEOrbfNi2bjVCKgdPBSoP8c
Ri2f/8ZartnvVEXNh468AQgRPVXcQuLejvOyRJXctkVBXc/PYjZMJGda2qe+NNrd
WA4fWyrFZC321KKl3npicT2yyRv/Bsq7FlMcLVQ1jAAtSFk0l47LBGupTzb9YwYd
oYw3ISpsX3alf8NThcRqEbmk6MWKkNbBaFZEntliSZAIOKe29ts1ndZtoM5Y4y0N
ZPz3bQEaujd1RlHYmKWnc2uKCxW0lyZmtllBybg8KXXfDpDRC1Of9FPPdSz14ONW
OH0XwCjQjOkvDOVa1BOuHOJBDLrVNCqDXo3em4kxClR02xo19J7YpJmnA9YHjZbP
RUcDHUzPNgbNU0gNxqqwE+rqd0K5+tvYNhgPOJpCHYKAQE7eNVRI9KMIzzspJQSg
RtVLBiDtFfpsITnjN54w5frA6XKp32n/v2cfemkV+ms7xMt2WdPoQoMqDqPS5PYy
Cs7EiPreDM5vNYCzpE2yjKfaDRLbQPglCnujtMZFJmYR4pHnxagCl8/R/kH8Dfev
PDBuFRF/rdoUKaI1OZ28AhPMCTBm0h+vaRlkKab4yU1fnxWuLG2Gh4cVB0fWFTuR
6rBZkEfFTVonu007uQtFhlWgNu1QRe+PfzszXRDvpjLJuD1qlkKIDAzIAn+l0G6A
+k7mZibiDOh19r0mHMnAtRJx1XAW1lDcu5h2fWIvo4FEUW3Wx8A/BV3XTROU2Lf5
LPPIOd+I/W6cCOIMSVGK+SgP4Fau98rDtTWMklPW6RnW0mqKavONG5TzLG+U9Wb+
0YdILZ4+C81/liA9VgIk1zmDRlID/Zbk9BEqBWW8a1EZoA5Snjxr2ZIfAJqwtcuz
iG0HxK8e7dSq4iO2HttU9hFAj85aobEPwywd5kId9EB8vOlvk6s6csDpZ3nt3Z0C
zUkarRBmkcUM63+MUixIbxt65PbzYnBNml+WFOdEUty//05w3n/No2ZSMDplnyJj
seR0RR0uBqsxxlWuZSppbrqh4DoI5aniDQftKUp6G0fwN9KadBLtVS20hBeyRFEY
AT07usL/J9N5z/vgQdyPtApKNty7vhQXJoa8lEkC89pq3WPIvvylf/oornV6Ee6R
9s2cpdUJ5TFUQajINJU8DbvhJClM/XEaLt+EBXACmuuMAMwU1nKOy1ElQz2yNrp5
CCMM7WdiKrIAEaZqXYKT/GXnVHpyLD31yysHl27oNQINybYKkd2QdKiKxooO59Ef
BlAYikHxoCNI40EQfidAwWe95+Mtmv4PCslg0CDsfhvalYWt1zgNPqtmrfYUrOwa
wXkgOHjzylXIIJq/IYTToQZqVdgZRvBLsNJSjUWeMX0Wc3TSIEjlZ6ymBmB3Sf0g
LDn+0k45uXrdhj7Z0l7UtLNxMOYlxAWapPBQ7ojAlv7sfNhgLQ/q6E49u4d1W/CU
foXmzxgF7j2nXwGj69eIHX77jSaFtfr9Ur0t4xS/nEQGLcENXrs/fCcrVkCGNKP5
LsK+oYXM+UHKokepXOJxV59JTmhoVHrfYTAYgLvEbRm/UnL/5CbBjzTeou8xtqty
v9u04f1rsP7eYvkNa15Yx9X8/7EwSGovR6Gtbcvw/fOMhP0JHaSKrSfpMOOpnf2n
eenMCwqk0bOvzW/nHJZKro8DxLpox4/BQ6IKEmjvkgbhn7cMJX+4pLzyWRtaft1h
Emy8ZjomZalXoNLFRjAHreq/id++AFtUyvZEwSPjj+h9ZqZWLisEU1p7CC3dtHsy
JMvJe17B5r379RKZzK7N1PufSZ3qgolYQH0OIc9rp6K4uRDgNi2YoKTZaYLfGrSH
eQAegmaXNyaXokUOgIqysBcyc3Bb7T9U9eKbrj0D2p7EgorxQMJ7synvRef3SKLM
kdVV9b9BgZKIDMfm8uijQUcd4Nyqh9NSmzgY6vyY3SfgxIuvI9uj/4bpzW92wK+9
pO+Q3yW2PwPUCOaZM1wxDB2wMf4WyJKWEexF77Y3d0oy0WbDQUyGgUwS7W2lG37D
ZZNRRpEi8q7wz8JLwFQ8aOjDzEUXs/HYcueCy3YIJcyn14TTmaG3uwYqYZIV4pu6
43mRQ4Y2F6mka9qzeRnkpCOSVzLjbW1E1r4LXpU9qshhfiUTZmI7VWXyYrInqsj9
CB8ePGy6uwAijVXlDHfaRCjNxGyE2IHHQb3ygaZ+h903xYngfp4Qm2uFlIA3xL5V
RWScTIRPGEFSdxnff1IQu6/iC9NUZlaKKBRE5KF8W1XXtVAqdRSIUoZEswJJfY5p
9OwUMRohtagjDpZGWAEQkggTYftyvs0N7XPCL9httvJ6SlEtT11/1J7lWi8MoDcx
QHir3ht65amdzk0E4M49T1lWJS693bJ7Y+IXeH10+TDI5qrReKOfdK+2V/INCoTc
+2Sy9pzQ9eSD8mQ8zrTbMhi3SFJ73HZs/1WU8Cpb+M1tCpZsakMMhug/IQzJlVfy
BvuIpBGLC4Q+gjlx/dmoog+HFzR9qpFPWqrHuWgf3ghMy1D02SATRq+IHZi5EzKE
DxyGy6GzGLFFpxn41l+FXp9w4GJ/tJHZH92V4hwgM52VrxyHIjpLTY9UBRwteJle
LpLRH8hI/xyYqB4SItSRWMOgXoECr9kIKHLlljUEX4wmILiu9txnis3+OzhJeZ46
3uq4nziC/5GNzRCQVlRxoUODBTCncYfnNIZXK/rDvj0XhH8Mw7YF/SMKfGvyqImi
yKdBetJs06UbEFvgPMM5ASY/fzvB37Jg3PFAbHpWg0zR2FViHOnQomkxs4cqqZTl
oCNp10uEcAguGYr4snssySkCfJKJe9ocMtshdLt4DJzS3nrXjTTtdQOWUQwmkSOb
xaZUhFJEOmG7QLFOpMR8cMMLXwWpnme6I5WAWPHFkuVrF3kAfsNl6Yu65Jluca0Z
Pm6od6z7Sn9/fFer6A7+3+nk5ShMN7zU6wtIYgLBA0fC4Wn7nCZdsALjEBopd5WC
CifwVDXzw4Yn0T8JEnRKfvcwKyyMPfN97G4bNKWY1TFQ9qaBr6T2fuPTr4CyI98C
FfGluCWNQ9jVcAkCD92pVdvJJNxeI8myrVxSZOS+afsi4Kb/bnhuksbpR+vfqjEa
VCAIF/015ymzAikUrHXGFqoEFuYd/2+Vtp47nCeAtFfZfpvLaZIQyMBX9LOEDB/d
EILqGzSMVSnV6jgWdrXHVwV55ID25lr0MW/L0QTV8hpwLAiFB11ZoPfOxFetRgU/
HhzqaPxmBjZH/OnLgQ1RJXLH8QAEMGJl9Xw1bJClCIxNo4NRij59qpU3DH1Qgf7i
ry4lXdumrc3pdkvtOVzyoXWJMf63AUwTiwbYyABZs88I3YNd4nIoY1+NkD3a3GKO
prinrQgXP0OecMtLKOSDZrKOa1NzFVvTvBJNlNe4EfH/OEdCRMitSHndGHm6pyDi
67BfbBaPL7lg7pfeZz53FItqGWDBh9y0SSP8vFUYDxkkwUV3qqY7uXzG0XpE7ZCy
XY401EB1D6DHIrMitZ4ag/413EMRc/unUyjf1wgYmFCNytsRlcc9FmSmzVCQuWgh
sfh4yPuPubKPE+hLnt1ysQHL6gnDapJeXp9XUsvQkeq/tn9FV0ChF/Odxrp2GmG1
YCTcFxrn7tCwewdSPV7zjuE8BkK7Nf+c89ZYSiuVsOKpFjdqIk1f09OTeiwzxcNT
0S+/xqgu33tLKRSI/7x1hzkGWeY1ABu8+HL0R9zexTnny4mZLr5jISQvoQWM/YlO
c4fO/3bJbp715+dZ5WSeW013XZ35N54NhMBLOEFoyyIi8coDufjuQQYp9LUQffA8
9NTWBCPDVFb5Vc4StiJAfq9RE4rtjD1XShmv+9CpaBvVUhvvY9NiOpA/8h7sTAUP
cZjH9qZlFVqAstXIrSmsis+sQIOep8RyNwIRwOlcFkeLOFZ1O6oRXa0Y8Aod1aNR
pC//XJmumjxJw3HdYNY7FrLO9SVKM0nR7N05IFDnWtEbLMkEEqMdXHyou3iojXWw
dSd5nf/VGqWPLtrqHMZRrTsGZfyn2QgRtqPjh2SNCzMMPEspW/KuYaCTtaZ/UMjS
t5f7yfSnHeD8zhvwFA96h7t76H9UlnpEiYErnKx/pGmCwP+lDw959muZY1BIQYKz
eXVBYno6o/UiRbGHKZEmFy8vfXB7IU5ocylfmbHIX7vtWndyRquhjFY3VrYOFHzD
XsVz5ixws3FJpbxHD0mJwUDMnXszGayNlsVmZvBcFJo7ggkHn/yjhvTlSq0+lTf6
4y8f/7vlq7JT7uSS75uPg2xeYiWZnKBHz/KGQQlz/SWIYG/zjFwTnSlUudfY8kAo
yI6c8ODuns/D9rZGUMx2lrH3XJvnzCHK3H1qCvIPBXi8FhoD/6veW6v2iOxAv8FV
meEHiE6CKE05dspoBvJgQomQOZ2IeugYe3af54U3fiWl7WKB5x+4NtEwpIM6OK3W
+Pd/zZ1sN+2NjLpLqVyx1OL2xBMo/cdXLQ98+kOuvulgCzSu0oTyJYTScS6nfdx/
zQZdT15+TeSoxs3Lu2qO8XveVnP13HMNWDb+PNiP/U8hmw7nEamsKwBjLGkhTIUU
k/Q97BmxmOBRxPhaini0iwz+AhmhlUMQ6oiXp6YAr8oq2uqiMvc0CvLcffbTgph6
TBoDe6896q5cflPAYO9IQiDndsOxv1Y8IgNzdrP+9yF3Xu1p2lXl12/GHVPMvPb+
OhF/F3me3QGbV9b6py9Obh2dBAWDMwHOSeOJ90Uy6WX0vi6Wh54/g4txVZIUdfpu
w4QZo1u6uZtuzdR4AXNexn3QL13j3Ac8VkKLL7+eM5P+car7XPG8nYVIZJDojYEK
cvbkR26zwzkaMsm3/woOjvicR2GxAUVFtGQM+fB1oA1yh5vvlp74hRPMfOvLXK8N
FH37TIVEQN2V2GZc1KA7422vnq+mNpQ0JkF5reOiJytIFmAhisdjKGX8nQKSr+MV
C7miw8YF8UYGWTIh8ir8DzS8RW5zAf2EOOV6zmkLxel836YnZp4UxjeHjFo17Wam
cANp3mm9g/cz1luQnQapExFnIvna0NABgY4Xg5Uwgv/Sv3gaN3XgJJJgxrYyxQUv
H2k82S3c+YPNIImvjDPY929bwp5xJuyElSWG4wD5NnI2Iizx4Zq9bm9e+LIbd+Sw
vHMAfbn3VZmpC5wni7IADewj4Y+PDal8/OfHmt4ZlyTYeNZscKgeVhRVukFoABiH
7na+YFrw1DyDrcSHu+fFXCrATfdoS1ANz2aTSsG3xGrQbHAtMbxtBaH92n7c8ZQn
GWG6pz9rb5KoakDy+gZ4ij0gjX2/H1LgzsfeA+heDkwpXiZ9ZXZFq71bWETZbn16
z1EIiX1Y9CfIOXbSXIzROt1aPEbMvFlgkEfMCQtWMAQ/ebYBAcp32dXjKXqDvvDN
CgJj2QYiMmjEnNVo4tgR0lSadq6KERTR1k8f+Mu5pYkqeM3bUv5GXt2MZKnZt/a9
PJfhv0s6Gi62fJ0gjTSbP87auPV3Wl77N1dG1OiXXFNvRecuYdKIYlXKQJxipXRS
hPousUW2lo91a/tKhb75EFsv1fdqaWuIeIK4c00Um7GBBT9p5fcAi2YDXYnt7gua
F/mJ5drhytiMQDgc+3HOBu7RAOSi4de6WCsUwPEzmMEvTouMXJpwJzfTuBxMGH5/
YJz02B4Zd8h40hVDzim4lP4SwiywS70614CV1O3ZwxMAY+Ioe2Z2q+zLGNj9VwpL
icZY8XA2c35O9YM+NLtlmXmGmOUf8Q/b7QuK0ndbQ1MMvlgsifqnHQlNTTDZWJ7A
3o/hAHa2yprs9Jnjw40PbGEmUOeRLnho66FFu0PNxLb/lunAdZ6DXo1u39JYGk5u
1hfTSHhLeN/lCQvloyKMbw2PNNfCRLdpn0s2S/0zI+di8qmoILhoj3j+xrIryxoV
SOQ6D39ZOpbT9GVQtx7FHfQwKZA3HUmc4buE0v1tHMfTjfSbB8SmZySaImPSSL8J
TqoK7lpP9ZHxdgrrKhM+7dvAj1HMF0dI7SM7g0ELExsc7Mi1dIHNgvD34d+D0cVJ
TmbiAujd2+MAkMIEq5dtQQ54P1iwG5JSrBie6rR4ZXKdNnRvXJYTGThiZoy6yPaa
/bTEEwhng0/Iyf2DSIVAikVA1aE4/ZI608gK91/QnMEKotDq3inLaShcE88ijj0M
FvkICOfYFm0SKMm8nysF/W2ci3g1Tp/hDJE24fnbpxoPSx0zeci+J8O7F+UfiXEF
vH1T07K0rOvfJ2A4BfUCNEEv0EAxA8TlVfhF1+cQNFKNVdn7BCwfTp9/bjd9p2d7
hDsB6APuS0q5v/nFx57LFuVID978nSD7OfTFjx8REfURywHMTzjPKtAVFeNSQw6x
3O32t5cTxhCBCS3SEdEuo1YcbQBAbwp4ujZfvvvCsxnkmSpKsGHzgUU3ee6nPXKE
O9lgfQTkg/+mdG1FuIcEAc1Il7o72TCxxC5WESBSRRm7aj4xLOHX2wCdk99SkZRZ
J8Rfw6zlcYul5W5ct8aT2RsuIPAI7rwh0dRs+7ztBHJGA4kbWzCp4mR4GpTw7exV
RXhqoCqchAuuClfnhWs6bcAOipZulvA+M2JKjAxB6DJGDDLS6GLFwxnte5dpuCAH
J96iFhMWJtCBeOASAn2QxxvvxagPbBqByR5mtC8cNvq8PRkaPzsbBnikZ1VGJLPi
Vk1kqlDzrZB9Kp/wgKOgN9g2zr97qy+ChKgP8mJ2UijtRJJsVyvkj4rgKlls0/FS
4PvOawTMjHqEy1vFT79F7PxNZ8fPI8jF7JhmetQpGnW584t6fVi0XYq6rnduQHvJ
LksGicNX7k4BNp5WTtuYZLgh9uPe05jLz/6/SjByUFvCBtEsenCVpvwqHuyCAjAb
tlJ4e6p8oTCne5hrO/vbJLdT3Q/F9qB545KM/58cRCWOxLFt5BN28Zyq4StqC87r
aQ9TA48DmAVAvZjOgl5Gyt14u47iZg2x/5+x6wDrVqhhad3hZxI/66ugZ+lvpklP
A66H/Lq9CLcauTk6ioyQvOsTmLydFgtq8wgVgxDgea7xFhuKTmVSXN8BBeRcrznb
OKcV3LMlx/O0FhOPOQ46y4u/eMtSzhihuQacW86xh/SbW+z5gbnaTTLlpmh0025Z
0N6EqbxJjWl4yaDPxp/rTMG90j8xRDTztka/dXVXl+a24ya7IYYFEa5tHi+xYKvL
sgxNitGRoSzRN4l2+D7/9dkDUuu63A3ZRAL/d6+KZWYgWr6TxJRHyNgfB6+/aOOQ
v9l2gcwUVd03KLvn20ffvTjFfhcPn19fp1jrevVOduPxOKigdlYz8z1P/dvWr55/
NALtoenvKUsw3CTkUfNqxyYEpmPCbjGxqUmvVHgnfnw5r8iK34u4KxvEbbAHGBjF
QWSE5EcA6wzCLWmtmyUy0e9/cTWWA/j9pA1n/iw09PlVxRkT8NtBlkTUGn0wOKx/
uXav1JjJvQY0svis2UhDIbUuY5uEJv38fGX+PssiwFuQ6JqXNQ6yj0FRSMKUdzDF
PJ1e+LvWxZgLG6l+Gtsx6XRkO+cn8vWMGSRE2/TipBS/lt+kLn5JtVPq9sVFklXn
9M8hxBcsY8CmKbXIFLAnGhyk9RLRTG34bCatoHdi7+9XTeoGAbfYZhQEy+754tln
1lL8J4McJbQnQdTCdI/KkOhZwMBGouuDMW/REmXM7ibr4tN5JPxi9IpANgP0TAXg
OrHSCVne3dNmY1A1F0XmHczkZbh/2Hk9drAYRCke9nYfvDYdOcSyW/gOdMYK52uY
ktgFFDgpSEVbJgWZB/vbG4fwnx7QvO4D70mIPOwNZFPo0JN6KFm9Iyoe9n3Hh9HH
yPBWSMhkC0uhYezaq5krMvFKofEg8TWUu/QjU7fTL+O/0Mlz5HBqfvsM/CZgIyal
V9C/dHXFDkYXpG0CsylG3fc+u3X+p+EBSXEPUDxKMgCE0XBnE31ygGkRyqOT8/A1
44VBafSCovIpFQzqQK5MDUxf5C1i5srBzXB5BQzrLL59WFJW0o1smn+zCugbq6+t
y2EYXNwVoKFW1VLPcP2aI/QwH1SChAlVY5iVSqbDDexhcynPlZv2WFR75EZvll7T
tPzfTyBEgvd47OYc+iGrYOqTYeyCFJPTBoa4swKqF9LGJwSv2dmzSi1WSqnsZ9Lr
zfS9WrpSWLPFeFkecU0J3RQjVVGOgd5+pWH+5j0yMZhwude0HmFU7K00sPibWqR4
ra/We9qtYCcpfjmbFGEqcp+nk1l1Fh3R148FqGIbTERuIZCLLZjzYxrrbYbCWiqh
MSHvoQNsE7hqIgVb9YzjHtIN9u//T7uzlM9RRKJ15JaAqGdS0prOgQYRLH4JCFZi
w2szWfQWXCte746LVuerDrC6RH5uxFVCcZGN2rPLezZGDEcu/ta8iT0TCpCuxE8y
XIc4YpkJ01Q9MpdM1xKJVzu0QuSx3eYayPlNRXsc6x8cjftRVrujdYmeEQU6DCb/
jT58sEHbDzaNAAneuv1zuZrIDeg8vRHDnL+TMsmamn2whV7O3DIOcjQ/62c5TfFt
Wf405sugZGrXnMaLD/G6OAath7v4+F9FyzI9QcNSSj2YhnFoHc40QP9Kbt3DxI7x
Qu2Kba7kN51zAOm1fy4X4IgrBxPF/+lin52aT+WQmthdQNJZqfMIW2utAlzdaPsu
2Egcr5kfZgsmXC4lLM8o9wCBDaObGMT/O+i/l7wZ47rQ+AjIEpWuSMV+FGS4carZ
SAp4uM9UbOYDsM/R58h3hqRdDvOucXxrqp0AP1nKZcmOJGSxb2dcekcbgE7nGITg
G0rnIeNIJy9ZSkxrtyxJGIYVmjsn9LzknAvcx2EXiXt9CChcoTDhQz9sn9GQFdbS
Th0CGssCvnHpAiNOyVlhoZcLeMzrg9YzKfQg3b0kkGdf7Is8DKDNNrFB5qYOWYaC
6jqhpzIQPXWzDVP4ccFVlkIOGWtqVV5H9A1QuzcHUBlCwoaqegYKm1bz0vlZPgD3
o4ZfFjvhTxgX4wilejz51aD6W5X31Oc7KVlrcQ68l9QdLpLS0wZ24hODi9XoYVlw
Iys9spFJZ5uiZ4qIYpPaqj85pRFr/tIXHAgMUhWdcdsDpBCGO0Jypa/MICnMzHyn
3qewiceNxXUi2smB2OYpzZscBiB4eM49d8jIcpTKvrASPlvXj+am12SrjGuwHAIr
hQj4/4EDkiCaHg+iwFXpUF/qQ76UMfd9/sEKnwNc/Y5Ne3r4zkOloncV2kGb/q/Q
8PLwfMtuIqFS8cfnkdjVAyhvVXTm24tDQMhbDRCcC7jMDgwYEx43GUu2AufeOEN0
+icUYSH5QN/fLoTRfcBM9p9qlHeIT5sjh0the7fPFvEf9v7wCLFEKJpjvgF+JlTu
2Ee0UlCNk4cbsDLEiUf9MFp7ZRkH0RiM7Mrzu0oQuEMH7d55fw2kZVd5GMH61DdR
5+ko22FRSg14tIKeq18C2sBk45m/c4nNmrWyHSC6CQaicDqTkn1no4v6MgmBxCkx
lX+4maqZR4FRtX+9IHWEhC0VFS6lOEQFuu7lzV4Nm20hI9vmnTazMz32AOk1o/VJ
M6LPO65MjEqdus0o6jT+VoyZ6x/r8S9gNDbq/9MgVL1CfpfxehyS77/tN14BMBVS
OpNPnn3vcGIG/bv6ADtOg0IugNRqDnkHpxG4Ry9z8sehL7JhbYPPmfo9EXNowUM8
p2EDJdmA0RpkmqkPv0If4CTf3EJYbNhAhVk4YutUDYQvEKNMu1chW9Zi5R0HCgNI
X8ZcasoiNVlSHKBhUMce1Va4NhGEyVzzTCIawweQbmKaZwiu/Zh2dJWZ0/V9a65P
Tldl1prBgAH1QWGTifQoASJXb/YUAhijJaetZRBXjYsJI4+TOBCv3oegpwU7hlR9
UShddJItLubZcFAVsqCNlq0/vYm/H48DOzL6+YpFk1FHCvSHJWLKF1yt+kuAIG3K
ZhEFiJx5ix0DuQgvoZEiM72Tajj4LYoCNQtx57qEB6Oap5YKXCbVpZ80oIB7P20w
60cgNuN+jWM3HHJKR+oQ7P2zgmqjnWp9zFWmK/UyGW+yDp/ItIceRNkgN08fuFtt
PH2QWAus/GhiFKgDPGmN9NecjT8MwnEkd+DwvbQ3BRZdlkRDFvBYDdAEUZSCUvL9
rFlWLcjeQZ4CysLIYMJeZt2KnyJ9Zw3d4EUsTYfU22XXSpby97TuQaQTukVCsezS
aRDMmFmmOakL11LZu9b/P1phX/ZBoa072IJjpumr/Yp2MfonAZe/8ptOiFuAVY5/
5h2hFUKKzUC1L3lCLI+wK5u340I/L90GTwcJmbk8DobE2pw665N9i9SEsQakzwC3
FJxoXiHZPw8Su6715IBHo7F/Eu4rPaPQj4Ybd2OUkj5s9LGS9oJJnm8ATLdZBW5l
G44jzunFb6zyWG/BMMg/ezVFPFrZ7Rk6wSv35JIeHDDTGV3+aZ0CiqpVTskmParI
GBw5kCMy/QyxRtZfSPlRPK99KiIxQEfnFl8IpUed0rLM++JVGHWpeUsS4C6PQx7M
c5dFCDI1ssHNtzA6Nij8WD+kmFKdlJzIq274rUN49N+V3mTmO4dmWXAH6V0r/UeK
ROn9Vy/91JTpbmmGi/l/mt8RYCPWzdbOyCxF/TplViwW/wyo60DhkAOwx1HoZa2z
q8hxq5C44tPW9hlUsYfreu8qGVSYVcu7gEg/V+2mlWJgWFS0HpCuNY/NCxKghjyM
BXgNF8z0XOK3xlaCoeBGxj3QrMzN9GlHh8vLNLi6elXYLWPe6/MG6rpu+MYWBes8
0qEzrqGPd6DwSGStf1F14aydyfbyZOwqRfccVuD+Mj8VplhnjN18e9mDezjAak3D
ldSgVO0uJR5OXjIblPCCNfpW2m5M4y19/aW+VC/UlAMOgzNZePZ/5pAJTOkyNQ59
50V3nPyCQqLh39sPTGimQRW0rw//YiJOw0U6VcYf2Ew9eOHDbfjnSZ1jX96iLvdF
elnzLZabveI5WvuH9t4UZL6kq7r4N+4UZ9IamLNHzpRtPoi10qRNLRzQpjvHD9dF
reUQEpSTRrV1ZDWr4+UhRXx0asx1TLdwlFoZjOa1+FEC9+vow6zk3qVv4u8Xn6Iq
Xnp1tgo+f7HYK2WK7IfCZ/Yk5T0xQJZpctWU6xrs8qfWrYszRtwmLNf3Hf0czF9M
a+qtFI2s2uv4JYN4LSzq6XMA0qmAK970DB7oVQygIf0kFsCX7W4X8dBwpMS6Rggs
pzJbplvNG4xxPOeXyRj4w1dmtMvrRpLewPEZ4SrI6tFMLdvGcQZgXcV73iWtOhRl
MY72tvCnqdr1plKriA/h9XNs7BoeYRPAkU4W0AuVx2KgXGYRdozyoSbQ5zT9q6OL
NQFxwJNtMUwfqnftvFAmEtCpVBhAF3XtPk4ROVC4EY+j9RUemTwbix4Wfz/3Q+TF
E7TgdIJgwu9MZBaY7skEY2p1j2PDsQZftJUpjV1hrQz3RiwUm1h1jRYokk/iMrSb
yNqzCedxZMIXdRXZ+Q79AChsFe2d3w0A7cZ/r+y/uVUblGa8LZxzTLizXvbH0J8/
ri5wlAsONFZl0EtIAHx5MoCxKMzEJnAbNGKFonUzDL2c1i72A3OX4n8G6d2lCBup
QaFy8nxIHSFjyCX5vrJ3LbMukJJXjTS7zaX4oyA2a1+1YGAF0b4r3afkqC5pcDiw
9+BnuNJrOE0y51Pis24GEq98JULkh9uTCFzrL7Okpz4kh/wj+hj+Utk4jr1vUpjt
BXg0TN4au6B+YHXTDdQqMUjHDVJAfzp5od81EPwaC4YB4vaKsM19ayYZ/K+h0/3O
0AkwftmUPuIVQwKrdDiIQ7MFlXyRhSVYfzOnVZDtkt/YBDqBqR8l3c2Uqkt3KAYg
OyubLpli5bj5cn27pLCIqRIZJjXOzhUE+yUmek3x0uPzq0606MemEbENMYUVVR9w
ozGGS6yZMB3Kg5KG9Wq+CdDSAx9HlTZwnjnVidJUurYPw0wyKtA9N9y0GKKdJcW3
6pZQwJ3ONZANPfvnU5jOxXRs4eIt1wCz/Ca4S+y5lLFkOKOahpF20PHQ7pwKf3dz
XH4luM/UwnYgiw+9lzzeolUS1BdBW/NRQAGR2//4Vx/pkqS7tsHfI5cbIcdbPK4u
N8mB/uQboRIopvfKSgFkM8GzlsJdeSNFofcniuFuTUgFndS89LGdJSl+HFyCJBi0
hJJtEMurg+GfELNucXp4ZsO84xO6y62NCFSKYQ1Fs0Bn1E+SO+EqtWAnmvqHvwhM
wVm/uaDyWhrzUBLem/ZbcJpz7Zrn87Z+75K+nBdxm5r9md5PQYPNIjmwspB1E2uG
oV59Tp63OlYNtJB1+G7sjNBIeYn0DndTnsz8off+BKKUuriZRTxzJsRO7gKpV9bb
jJelIsPgOdqN9v+YKicx6S6YBkbvaQoLNxkEu63vQiw7vyxz6sk+aMrk8Z2g5MNp
7PpRXt5UzE0CtBDIWJzruiakxbb5YcXNAaa3VDW3lstKboRC7e6D4kSpnZFzTen6
XfrZrqo4/lfKvQAVe2TQUCEYIyCDiCP03f+ZsdPNSDHAUkb9vE2STvHqWSoyzZtw
MzNKC6M5kvCh6J8zjwrU4VbrkN/dmDB4hxGOolPjiBVQbWi7+ECzTkKLfP/j8ZYD
f1QFKL88gBG7izZ8vRSZCKw5C6XIDQ/pfSo6TeB19M1yB+Sec/1E1qZqbMQC22xB
x7f/bzTJnUkd0/ffXjX9xKko3/foe+UcOi3oxT3AfQ3NRAgQEshBHW6O6Sh9tHx+
UnLDqYQ7s5xhgw1KAlkZqqZhPH2FQYwkJYJFECTKzA0vKn5GfIgSaO4GEob322r0
uxSCRiVBwyxnm1lg8lxlrFN+N3svw596282rTF0EoY+8MH/splYlyb04SVA7SpjE
7dcGX0dRb5CVRb4fWmUSkeIzIC3w3qi0Jrq//bPLUDmXEjwLfi3wX6zuxRwrwONq
dCJwQlUA3bQdS/ymXVykBJKvvJk5d8mhgCDPJ2v1U0kjOBZKhdWMNhbG+Fq04uJO
GOsmrrbTL+DRSs5YOSzCd019sHRWXYJABNwz3GJIzpZWm2yYdgyipVCQdjH99wlB
FKWng0DswYRkOxyFPnLRvFOMwa9FHvuf5d/4KZh+6dnDPm9++KXpkySCsWu3ud+o
s/exs82tcl6SKFDwjj8QLQt7ruvfsEGdOn9R4lkxp7iSiPI+/5DKqbMc0NdJtA1i
m1OuX/wCCTLEJMYX9UilIGafV/m6zskmMdqehbF7Xl88F0Wa9qCnUIWMYBjXeltz
+MCvcunpHVdOgSNvfPVuvQoM7BMUMAk63kXPnFjCzlhOlKnxdQGxdLvLfgzFTQvy
mpgttztGlb6cNXe9AZH2MXW0exWwSXBgOvjcIppttwAuV9w8BBXxlakKVXzGh8OT
ShxsJCPfy6v8+r3WSUhe7dDjnspGBO2Qz7/cv91fD0uCRrBjl6RM0QvN6yVmvLlX
uoSWRbONyHhOavO8j4u5Frc82DPUuD/eGufFM9tptAz1QslELFvSMHQCwe3HFDun
6SkKoz6JGdmcq5lnt7dwAQQm0FDwhHzpg4oGEYJYIYPxlzJiSqED9fH5znrwfAZF
Czt9lxZU3VC+44iLay38J/D/NV2zUOJ6zkyUFrQChRBonv7wM1t/7Z1UyXt4cHji
Mm+tmuuuixNHteQM+YADGFA/HjQ0WdqerOuF57CvqROZM5OkGYtacjP1RAHxYe8O
6snOG9A8DS8Sp4V0tKypAQcIbfq9DA3WWRYPIN53sSnqWXdshsrkHqFT22CQcn3z
Eb8HRlBajUEcVuL1KFJ6+njZMAYqYFE9KS8Zg63J/1Wg8iafQPEKW+0ujdMMCJ+L
NETCxsWK1o4bsaE2EfihuV/2RoBCxDA2pYwAfiuu7k6AKZd1UwcWcMQdiP40ftcn
65xtzVlJNYVQsQPUdNShGuHMNednuDHUJeTdB6qByFoXjfFJ2ftDbIVm62S/MTby
Ogs1sUvN+Cgs9zOdos3PFMUnUTr0GQtK2ZFzIIGQ3gJFdAmw7KHPvO7JnRQIxUjm
3wC2LQ7iw7hy2CdRBTm3RUui8BF2Qx2SzubTqghgBzA7dA63OitsSH2sMw+2FNXk
tdZw900/dnwaHXkfvWJ2zLBbFjbDGxXqmezIz9X42SGT3H/6b3T/S3xnE7LKUWLJ
pP79Ym2oO5Gm/yIH5Jo0/e0zVQpOGIW8m9jVObH7JHqIn7pqP/JScoUZUr2b99a1
hNgCVJxNwgoNvw7BasgNeK7/GdMzj3dgGuqNqRT+9wNwmAswq841O7LEG9AgYpT/
AbTaJ3gQYG/s03J/lqqSNNZvNcczZRObsdn5x4QirlhAbziXzGzh6hooC8i33W8T
Btkc372LEF06Ulv6LFtCBRg430rsWGOi6NiO1GkJFBq5NlB0apyLdS9jwC4VpqPq
11BKZSmMO9UW74yT1rmM8h6ipZp3pmZQquH7nPFMnI6pncqc+duSY5NsSfEKgPTk
utw219RdJsCqyk0XKwvDC80x94D+bP6NFCa/5QYPWCyA0LOucyJOKtvklIbijuAb
rG9RTUI/Oc2dKfBUK7fMmwLsWnc/f1Sy/Df9rbX1BxWMhpFFpfy/Al5fAX8WA5kN
1E3OH7zayXq5FvR0aCmtYhHW81Le2lEs8WnrMQeBpv137kHR6udqLBtNrxyjQFOY
nUfUtW3ObF5qPFq14xiGuN7I+A8i0pVhY37BpSiagZocu7JDorCI2OKOxPARBhoE
kt+N4pnrIOlrwlZxwisDi57xWOL4hwNxOfok28D1KUFPZ3fKdj4FxiJTM1PoHJQ0
d8P64HIRSASV45TKQH+HhLq8zRlp1ZCJr+w9t5FT4BF/wUgto9fica+nolN1J9BK
0pvj5kC5nvzz+tzlB6MJTDrwjHgIxhcsvqtOnbjbQqo0vWzenGKhNqIYyaQnfd2Q
xTxnBVYzhIUn26IbiE7sYQRKB7W/nOReBGbyIz3sMmhyrLT90AE/x5mYckaCWhnG
WAvjdb2RoUXtTsZTO/GbaPaLKHanDt81aBpn6EbXHwwmUkkIRk7KeHeN9caF09TV
qSGzhPCycUf4SHML1Tbcne/RE66EuTjGqo8G5m/ZA1gn5XekYEd3yh5Ak1k4JG/i
mmUOyCAdfhJLkj2wAagQ732XZ3SYhN8R0QWka7ZwNbE78OabJf4ick+DQArcC8Ii
oC0Jh0PPYjf8+WAF6jJCIAF6YRCU7uNXWZRnsSrsLUzgHnLUbGVE2F69vuOwPa4a
lcT26ch7EsphkItoDSTS7B/M9vIcV9jf5a6ki4RY2E3Y0Pu/4JXsEsv1tWAc3VLu
AQIHOJDyNTbJ1X4XrnuvaZ9UaNJlFwFE3uKUskxS/tXBLRbEbtfer05tPwv0X2Iz
Qju9P7mHwI0X0Q3wY0bgYos3Ggw70UbmJQS8irqTm88hTM0om4SzdIg/o2O9N4Q4
x/Q+zIKH3e0+Gtnyasji/iB3GCpBnFUBHswLxppnIHMTn/1wnUF3cI3Y9CVyrPsk
l4GOuWF7RsRvPhnhgG591+umjbHyw/ElC4v/pdhMeaKCfHAAOB3Rbp7BavNlxZ4P
jtenCYeXlEMbwc2eiPli9y7VJxdoBJexU3/Hr/1amTZ0AiUurFKIPXQm6ViwDDSk
AZOuvcEymCL3cpnVenrnpqXL91B8V7J0CeaqNcs1M0dire4jDkyUqcGX1fUnNAaQ
QUPhZ7xJCHzhI8iryRxUs3Y8N7TG12fYVviBUTnFWpK31ONR8DLm5HpeWiBETGPk
S1NWoWb3Dn0o+e2wuktxW5DWETJs3ss4yZgVDkyHC2BdwNelS05ws59tTbwbmbRO
iEeTQvNzL/l9YpIE5x6YniauIV3ldc3SPvncZnzPNrQx5n1wdGNy5881xfLBhoJZ
IKmeBG1FQDi84QK53jeLUcfS0hEyB3EmrNPxupbjjMFyTp5MGns6u7eHtJHXOp8z
ImC1R3Bh4oUeNwzqIyxXhPzQWA0++IAI2ATxsGnCxG9xDmX0Yf81xK9ZPRf7OhzV
ascGtb9gLtpkhE7K35vakRybKF9Ls9N2FkvbOlZdw/+9Jv1w0goKIIeltiWMAFD5
IOAOChRnMffr8TWSnyM8v+8WalozqZrHfwL2xRVBpeo67SQldnPRRTPHJ7OiNIKn
67qzZZaSQZBIV+rvllJg5BflVprLvfhhZRGaiNpeg8jzlCtcF8L6LIvoDK2pkbQx
K05xjKwRHlYVhz+tyfxfKVJ4q7qOyA6xIfM+on58A+WJ4sFkolPtHBj4Uf5G1/8t
3NGhM7ODomBzj8tRvcGPO8Wp6qIei3QAy1r1I7mZG6QFN96jWzqsULzV/1WtMa6g
ea2107UlQx2JH9saG8RiOznL3skO3xv1llrzPe8GRq228sLrvUMZnSvEaXwvNUe3
YnZ32ANlVifzV8blRH1YaT1Jd++6/P6r9H7BVAHyrJx/9IoCXgNtqqH6H3xQIibT
ztZj6MAgnr+uQqXUFs1ACtspbLwSkK1hHellt1SAIRlmcGEUp6rFC4AzOj3aIbTm
F0ePUQGLqhe9Ej3XDBeI/z6yMdpMcneeFP6ZU647sCoBWhFzC/NEwXK3YnH6/1JL
5cCXHIgWZwjI2Cf+ZsvlnK0Wb/nImEOif6bbwv+hR6ozUaaL2xTgfKlw7nMl97y/
BnGjMbJb0RAIjb+QE8XExChHHsBcR7hyGdnZ0I3htbubK2cuGkOnurbcyQIzVTnV
/5Z4h+m/TXMYla/scubXTcyiTEiUOQxa0JATXrsSAT6I0P1TFaTuP2gk3LLpCxjQ
d+th41D4m3vGAcNY0dWUXkeThF1WzsE5k+713odq1VeZMXXeb0s6pB+U57sQkuXG
mZ6cYm5CWFXpQHGHxrwfjP+++xVxyxLCBVa73DadZW33P6WYJ9Yat7G0+i6KzvbQ
H7vSX4ykbaYAKdoH14nA/2IK9HOpjwgRvvLvaeRYrPgA9yOY8EJMsBsgHOFco6GJ
gGdcypm1+hMVMTHHAtZvceIuYXocRZNaX30RLMUi8pC1lI8zmcvVH6HdudzjGOmI
XwZwpBXmrJJTz+5hXsK2zTB89CDxec4lWI53YER4cZZYJPM1SwOSVJ9Q1oeUsN0v
h2VsXp3YBvVBfmcjqih+rH+BXP9ZBm/1v+5VCRcMnR5k1j2pp1sz9/ANKGgujLpE
yM8UKTqJhv+bLOJg/KbrclPWadtokg98P8Hyi+qQ9ReAKb/edtd79I8onlj3oqbZ
UWsxvxzop0/mUfKO0ZRR2te+OI8N8/9qX2i8xCAnnbZLe3A/fEwePmboXSwcHEmK
7LGUQwCX9X7yoMWg25vhnKZZ/XHrR2DH8yvwTR4scFLSvv9xbByxfSl+os6maOix
tbEbFJqIwkReTv0x+SIZIK82WMd1w3fPfHP++KmOAuSLXZ5J7jUHouyPvHL1w3MX
s7j3UlqTeWOs+YZeH+sqze+h+e07UV8RJ1CqkBV20yEXyuS1P1bhiG9QefI2J+Un
gvxUSKnotPXDzVxrteJ6YM4Yl7a69adD6kFMjUvGKTFnyE6yiO3FYhh4TM12bxMN
gby+nhy39IRBX3LKHA4Tqk9LlBbStuBTG9UhI2imB33Lz7BhdJoKLLGf0drok2K3
jVjPyhI8kUiLNev3Nrq89bJoqYNL8ImwtsNpUZFlePZgledUA3t+IAFcEuU9ohy0
B8XLNJJ2fVsca0DpyDbLqVD2O2rApBvMsYNWkH7dpTgLE1u3NgJWC8G7Cmpp9smo
NY45MpUWSJfm/X1WCKxJZkZ0OysJ0gsOpFrPC/ulgC0C2/k7vNTsxGQ/ZsA0yZRz
p4xa3dms8Nx+eaMqCGQ3eLnt54cixH34sp4t4NXvt2Din1yWV6mit1JsLoDzQBpI
36QZ38I6EgFu2TgsdNyjmCQusJZYcpe/vt69otRXRGY62InQbP/VS8XdeFVivLlZ
5vhADKWaLznCnLMgrRBPStrwucYI0594YCqrPx/NvuSKl4tSrmcfPSK7FlyiItZL
P4mMS8HimuRnT0/EcE7CT3+UmcNmk3OV3ssL3oybSZ0IXgqD12a4nTh1C/82S18U
InxBGjhc2Ru+WPBqgWlDp679rgarG8nR/wst2oz/YQNJGn3WlWwouk6O5UdheGG0
9nQG7xQgtN1JLpGvSGFbkJh4s2oqDVBCEFadQNsqSX/L67Cvw3RfC3grqKvKqfT9
N/cP0O3S4WTP9Opw5aNpK3NHHGBEX7pmpG4oqu8Ft3/GIq/kVqKchr2OfrllsaX6
Vs8R5TkNIaqP97vDPH2eb9ihsAzs2xPzRibW+dewBbHlr4Wly9xKtLrmEmsArL0Z
qLBFrBKF6/2cAp/43HcyYDuCLctRm/LaS8ZaCL1WrkV8nh2VyS5sgSmxpk+aU9oQ
U62KRQB1v4SmSYbvcUtJ+0d6u8K8EzljygfbBp89dP0hOQXpROSCh5X5iKIGMsL5
EuS9O8ftTJrzTgGrtA5QvKG/gs2dejb7xKjzQ30YIpy7rWji2S7Arj5THmCFIF3+
FjrrZttfhqs8YmZ3Qwt87Je588rs1Y+pXtSX71pqw5WJWEpZKG/LU5vN0phavxsB
72OIxfH7gCB8iEkaI4O4VC+XMCKhdEpRq+/Gx777261FJOuvMqwOphXvhcW1vHLr
zv+fDqdOIxhBrGld15VXas/thI7weMAWUOwdsSbKRtBGBuidu4Fd2Md0Yf9EPTCx
xnoILQcRO41Za9L7/q+j/dnVJRc0485bmgWp4ciWYf1G98YTVq0Kb1AKwkqPbNQa
58kXfVVnUAD+0RPRxofogV1+vxhgIGoUI6VqSn+39Y3X6h9S5IBNIBlcnCu2cX4L
8to4tjRbVQMlfTgAxmmjiquCP392bVx3ibXQRh3ujov9PVVHOfPC5HDAmTal3SAe
w/eSigj3uGEZ17wuGY+lbVVPPMmpF57N6b8exY7b76l4ktKVmgdO3XwOr28b2wZR
iMkaSAEHA5skK0FXwJ94BbMp1WYeJkrAWI/62A7alHnAHTFIrWuyK1l2mFsWR6rp
Q/MdaYiS8fOy2pknDxcHqjRD8j90oZ/lixIdd/jSXEJ1Si4QVuXDYdRbXokbp69n
/xSCSvr2wwbX6Mi1jODgLIJ997UHtsByeRU2157WfmZ+UnE1k0oiHzSggRe3BCga
cO1Mn5/TaH08breAWBsJZgUyl28Sfk1Ywy/yrb7KPDHYS4PQ66taW64S6cleUeGi
24Cj1loLwMl3UZnIOaXbObS4QwFRhp/YsbOPHdTWTJ1JDtPx0KgDPumMHxeYyh4G
q3Z4xptpeTHNYmtysw2Alc9pj0NCi2IQU4mrD6Tl4y473X/yJ8tKjhNEirjDwm6r
1cNh2diZYPNJ8b79kyaEr2jAmm1NSPZGzbMaa6LIUREkOLkmNVFVZxFXunOIdQJt
g+/p67rc3mDuZsvjJZ5mv/xfdIypu5MIn9jSK/TmEZc+pNoRjzB143mAGal2WT7n
ZYA8BNOLcaOyQyemZnpsRL2z0hXjGf3LEW3ZrjpkAlOAFCkEErLtd/F2g056Pipu
q7VXVT8CogTh/LLpdOCh4MDrE3YOkBIAVvGpNMtbAiq3tIbRNGwZreoMKUSW8oZx
1nSN1yitqhKynBAxy4q77Nt4e28WbQXdeQJgd453Y7IDdImunY+xZs+X4V01SESr
tP7OqBrmy81UE0KMbo3lHJuij155nZYCP2oAtuH5YsfEmNXrMZv7qBhfP+Gs/HAR
807mC8DaHSRCzx1QV72pwFQb8dFVSlvkdZTYWgEAGcxa5jfeHs+lLyirRsHZXiy+
YY3xGiCkDWXBBODHRkl+wFGP28TznVaayCUWga8HI23+mGfYdK8DU8GgFukfPMwU
dkytXyPNbHnnSgrYL/++3W2PuzRE8a2SZNGEvcE/QJVEO5qh6bZFAxKhkmB9dHE/
GctiBScey1wYWOqzdi2MN+XJ/2HRNj2OGP/LOJi1Isb42bNfvjzfgH9vyOFp7AVj
jiT1GU4aNX9QEJhctXrMm2Y6u0jaskDpGqxIA848ZNbVPFySRXkCXokTsZhTrLAY
uvRHGN/3ft95UmNmQf00Lz+KObZF+eWvzq8SZIpe0zm/vopR/5zgr3T4EVuP0hoa
zFtSIQ27b9X9vTNTsit/O5t5XPTb00IvXops3bSbmyTScLZOp5eto23QQ2k/lXqs
WKRzowHfi1IsrR48/W0wKSDI+FlqfXPWeI3qB2YJdhRP2nQo8kbJ0gHyOb2DeJOb
lUJ/+PiycEfZ1vRTjPDPwThy4G0IZe/Y0w3CBF1di9Y5GT7gu+4THCD9uumr107d
ka6ZwUyKsTzMopJ959W9NI+RFsuiHRdl2B97GOkqVeAk95ReaO6pAfU2ve0VA3Kk
2QnYygRoFyoem5BucMw1Z6eupzaNRBjlnUaVPLzZHYo3I/LyJakEtieUrTCjNvmD
DtgopsvOnogtmroxr0zI6qHo06qO/brdWQJ4w55BXkg7VkG7fE3TLEXVNIlJLz5L
LhQ/HwlQwLeRjpJt74BNyOX50gE3niuCSGVpFV1WDwvKjuP2PhgtFrL0O5fca8o5
Lj6nn8iOitiwUaxWBEk1HC724/77LrFEM14tg7WDeOpedwwKAWgDlu6BzZqNLGt+
mnwDl00vTFCK7cYgcZ+z5MbY4MXoL2CoJD6VFe/S+T6Qx12QusrkoLRWwQP2e+n9
l1+hQjHLuZAkUHFVuYSmJ7va0MnPO2HVJZMYA8ElnbtCcGwYWhwx7YfygK/x0qT0
bRAfdv0rcf8d+4iGzpwJ183zubcsMnp47kBfaHU11J6pb77MO6DH8GLRRWaoBKBJ
hcfMSFAjk8TRfv03z0CCeAbe6jXEqF8qX9IjOJGCNhGZj9ZDzxkLzGZZ/81Zp0Ic
scoZtmiWZ7ODmHlBGfokGcDkbtAMX9ZBjbmfbZQy/kaSMlXBkJXplcQ0v1pRJmbl
9/YqM3t8BSOZVBMAx8rm1iZeu3cFrOrBEn2Ti37CeLaC+XtcWfoQ22QjIbaR5ACl
srgWWJZY/Hfp6e8KOmzIr1xn+06bAILTJBnfW64GvyaheAaYwWAYdEk1ksa2IjbT
fb2ks7zXjYlNVZplKu0GeQLnYPfRi2grwfT9l70U2PhdK2sNKahNW05fENdwwRb4
aeg/gAFBeZ6zsCocdYD8IFqMGHJ9HJ91/kOMwJHhEd9Dnveqol6uKoOfPpt9GwqG
mgzwsRQako5fSJqqQNde1x0qvacyi0sMQc6sagamvNgVKhnYdMbc4GVYxarTb8xE
Qz3e8UYt0wsmsCAUYn6QBkD7B9utustXhGh6QsO16rQph/MIqn8eQDDsUe7YsLnV
NFLiOhmPFIC6a7YTdKLXptQbiYqnWru2z5NfBkBVmK0kgqTZ+PHYnazLycy78Au+
vO1bHs6z6m+XuCkfgBwzJ3IdUNm3OhmxVdZa6ACT9VKvdqd1i/pE0uh9jfsdPnYP
NFrjmeHBvcQfyKZ74th49s3VlY/weL8vVbnQAZSqoq2ZKBpBWhqZmAxsbNKVTDet
Eg0xr4NwOMOiGRliGS2Mg6wLM3iKjFz7PjiHPGM8rutIHaSvkzs+DkxkqngMvXK8
krQOc8vsxCBXbARj89bhT4U/xeVaXQVxqbhmsIeQzvmJFSrDIl5TtkAtDVEkY3bx
lDL8V89Vxeq42vwT5hz2LnXz32pQVdQKocDEc+DGBa65s52u8t8Sc65Xazr5UjBm
MsJFTaFoQjP+j6hMWydxNw9UovPc5mRlfzFrHTVOS8JAOGgll+D1CKWGN5bKcTqJ
Ff1vnOEH5dUtJyvBCYHBY7po+FFJY8sJvHGVXN6TlZ2xTkPtXd1RZ98CZebBfRdc
d4Hvwc2/Oyyf/wONLwd1Vjl2sTHfogpGJJYbwxkxoIC0eap5R+fGN4fIqUpKm38c
U3lPy2axKw0umfO092Nojge5jlCvQmWbyyFTsF0VfvPLEwrJ++GZ1jQDWmPbVv6C
SgU41d0kXOJlVHFZ+imRwnyNeIIHAgWHe+ZshnhtG2lSPQjTYAZGabFTG4eXjXDZ
Vhdg/C+RF7qmFFfQdv4ekUKBsdz6UTtSsEismMKNe3t7WEuqIMn0bgAirrqlkI8x
b3Uc3/npv8GLt2L6XQ+Wtk5Z4TwU7h18pP4ZpHT6EXJugHMUEsc2LWZs8o8JoHlA
Lz8tgqEoJIzmMGu6z+dTAoXlSR/2R3k6UOqm4VEz0J5wPRFJ1x+7lDAxSBy96Ycu
obC502lqlKd/+sEKyUjiHS+SH0rs8B4E0JIpUX0VIILdIsmWczYvHMEYRsCl1eze
giy+7fxu3ccXHSI7r+rNCSf2GY79NavApz66pBk7TPOG5rKqrCOzbKtLsycZmhjI
jBKADe6u0949hBaIA189/pPjv9IodA9buuR2Oq+hgtLAgspUADw84oL7hdOQzXhW
nKlY6LuDdPjpycNK6qu4hM61f4JIDCUIoPop3CcUekhpy9M+K9lEW9xHupEELF3s
wH6zkX6VqMP/6JZlLm7shETBrGTntSutLssX8CmwUyreWKGeBf912ZuXNeC1XSO6
hcRARGB0Zw/mWEiF+d/Zo9EhvQ6vvqPoxd0BSTZ69EqtTUjc6+u/Gybab0NcX1k8
G36le18UoKOGEcKmaiNKlPBdhNDwJoefg24HnkyjLXp+yarivtmDrId2/E7t8PJ9
kNlpelgeUAOtrrJt51rX4N/eGvFHUwpztP9FTSfF5IMdmuoYqR02vre5hAmWY9m3
g2wqWzCpUb7eycx4v3+ht4cAB2thgXuL6ueyGOf5MJVi9TZtcmsssxhovS6ivJEJ
9vQH3VRQssdSNM0QIwObE6vcM1FNHqy4SGzKqhtDvWlMdkdxQITBxve/xfpLdJub
2WbcajOSnPb1xzE7F1zy5g4ZrsNeIhnCalEzAZ2Q2eAyfmbE6ay9C9giF0wo+Pa6
AVd/B8sinqQfbZdRTH56lxs+pbqt5jCrd9NK0Yr2zNo46ARGZ/vVNh86WylWvcf8
EUSUBEloR7a6Adaqi4OX/8nE6vgrBWAWIjEIFTeleyW9xIgLkqPH3no3BW6j/rtO
CQdSKyACw3V+eP8sgslXPOY3+mhhyhC54/eL/xbfVAh5M8sx5Sa9jPyzoTn7JQkJ
7JtF0p/oQgE5Acy5ZtXjwNGL7zAIfBaatKUINSMDVdULmsHb542tPuMX4QNK+VFA
rsXPSYahnfCO3UcR4/MT6NYWYasdbxGKlD3rx9GoeCjg4LicvUaOvQPBFbx9CtvQ
iPtnnxdnpsDw2J+KX0Dc/AqUaP1WjE1iohL9G0XKVb1p57YUV2HE1Le6Yfc9CAPO
xKp2WiTk3E89D+5ZAHoLvyMmJ5edhaSt8I6EKIvVlWIyV8w4/XB1eAEBWqo7ALFx
lotizDkvtdURO7BaqT5PawnVKVKaJn0uoEobd2YXFUXTIG2UxXS1aFq6ihKrtUzI
2cFA7H6SUq+t1JaQsRCGhotYtXX4oyvl12X97FyItd3J04/j8o65Ku0keiofLLTy
BQ+BjOM9aCM3PH2t508AxUlciXSN3TxnJ76yx6qWKzoxtiKobemitAB+ldXW9gP3
nWK/hcJKIkXn2Cd1A6hwhGkH0P87K9J4VDJLG8UCBtjbEF/fHhxTtYoMG01au30d
trGuaNbqjL8WTK+z0kdMhzVy7YLDtwOdvzmcnC2OoJwxxzUdMcTej/G/fb9nUjf9
hs2i73IlhEBBtrIiGOu8/dgj9cnVvda2uyJhwyafqXM1KHSByJHgXOxhiFvf3rZ8
r7rXdvPqsFcdacNiLXWSWd+kEz/3aWcVWhDhwP6tDEHZVLgIBHRC+yfganiy2fbq
m7lrzmsnAb+UUDRItPpcBvX+ngcCEla3MDf9t6dIY5VOkPZbLv77Rt1JyZ3B1HaI
+hs0saaKb3Ms0lQ6mFu6HYIJfYbMSKkfrIR7yBpD7fB1yZpsd3GpWJA5uzQ7ApmK
3KLLytVk5lQ++ykfJq+RvsCfRl8sSAnU6jU2mWyv71OnTYDsEDSuWcmqIV0VecY/
KrxmjP0R20r2MbtB+jQGdOvK0ApbIP6v559HzbQz8xWVLyozOOzt46AiVia2Qd0M
tznnXkCbFduGXJ86JY4aNWzHwdlveyXft8CfcIxHvYmwy29k86zswKGBsMboMMCX
hyxgApMnXvfWnFPQ5OfJnJBlMkMXGMNQJm0iBdXKym4X3Mli085jQNmBMURyn8xm
S3lUR+X667VMoYhQ+Wydbi0GpyzwaIGGPAqn0CR8cAmk+DvUJkw3KVPWrJzZuyA1
g7MPbM5z3sHkSpSFsC/wWczQs6qlrtQRaWu7AW+OYcFgq08I601ltUn7tOszqf7K
uXkEiHJcxzpVAEMsJUcXFH7RMaEx1ciiTNMWiPBsAousSk6hQRCUeuPxUlh4UTLJ
nBGKCCpGe4XiJD1Eil734XVjDrs5Qj6d7669NXNbtu7y/SdnI2wsdDvEE9zOnG1y
0l22vchwWxshm3CvLJ+yodgyMz0GUkrZEGktk5t8cQpw15iHwzicH5IXWYC9Tbhh
eNwT6JADFSKX0wGA3g93rPzZQNIsol2Quw+liQ7a+oJdlhw1Dz6ugbOpL/Amdoo+
F5r5gKnvbvhuXPnppG2YJShdK1DSEmfl/RXr8zwx7O6nY0P19MOZrKIpRcDSCxJT
OeNuj7Be3WyhXS2qMH6u91EJaFvl8LGsTU0aZedFHUssOuLoK4269JVeFNDdQdlS
lbA15rRHKCPzsJAJ96m1xqWaAEFI/fAnkenZYp9pMa1aZrBGWmqrWyBFD1eQ7Fj2
0GjxO6Qw/O1INHkLL0N6UWUZVtJ54p9Wz37BUeBPq+BaAOocDOEg0dPO9FYQ8Qof
CNLlkLcc9n5dPSC3jh/O2WmgUZLoPLfs3F2mce6u+zFygVUyMGU5XIIyW09m81Aa
IFHaWWkJZJMoEU6SfYox8jtc3Ck3vu1D7xjB9a8Q5T8hkonKArTglNku1NneLie5
SWDEOFv/Y0mtPEIulK0/nfNa5XNOSvjofRXFMT6YQ66/ZjETSLiwFFnCJeVgD5MM
UhA+lPEu5bkP1Qwh72lvapsvgmOR6qITcw2def0rMBa6TT1AtCKYx6pYsW0A3wyh
uTzBj4sul+n/RM52hQ93Q/NrT61weRnBGwiet0zWeG7b+ofV5somGEtStRApfk1d
Gx119S5fszSrFEpyb11Uvot3TdpYWD36MvYJcdvq0xEWw0yf09oL8faLafjbuxTo
UEJkC+p4QF0rAjGxpCfno9LB3lwW0Ag9SiweBAT68vREEd02NSaGUnCRNQeUFLva
XveIjy8cObSKX1EFxvma6IWqN6aaN9ASsAeEAlJGFEZt58SWAAZxs+dOGj9PvBbx
k5UmRBG6lPkt/9kADF6A2wXxlPvgQ/9voQ1mN4R17DAkLnH4thDu3zMzaoQw25UK
sK+5bABOfmJeasdyBUW3smXV4o2pUFD0fvmmgDtgK5ZBGVMyluwlngtt6Kf97YnB
kViBUoAbffpZbosemkvV4S4J/kYWuwCFobKRuIGx6c6UgEsMU+deXLGm+x/GDJTg
ca8zsPBJFwETLptUMBXF2kP39sr75K+KYfdrXz4cTFNmpCRdRrRzyTSiQx5wQcqJ
upTYsCzE4r4Kw7U9+dR8T8Z9jgPygGs8NHvgof78mg2/gzbvH5gxUY1YVaDtN+MR
mU4OAOmLAQwU70Oyf3a3BpSUCikxy7EjdHX27d7FrcEAVt4nf8Bo5dRm7roEDIR3
m+gL33G6FV1bgBh88iL/UBoXpf1N7xhxlPMryskUkF03ONf+zJysLBPGeRmQrJcm
f8ImLdXzDAb7f6dTjHTogk3uWZ6E4QcqpuNZ/bar2cu2buYw/VsMSSbVaLZEz6ZH
iqn71S9nRcf1fkdiSRt7qdpagkpWVOBLw00J9+BPjJQUaM1kouFHRxoOmCRmn3lw
T1Zja5yR0kuwUd/iPv5sarUADFHEX1Wh07XwJR3HKIvGbUVy6oV18Z53Ka6Ki4of
A04OUE+Z6IvvsrzZXxyeSgGOwJE0MG/AviiX20dsGyiOegdWjZFZPlPSzl+ZXWIM
4fvoaRf0jHrZBjr+Mf82P9bqmKHyJFmYFujar7+9sireG5bDdXRYF7gCmDlD/5zQ
LlQOKp9qEaCaEIMS6FDToXqfuv/u+zzf9zi2V1vG2xk8h3gpGFS6Yv36T3qPkOp0
zEXNlL4XV+PxClnWZEiu3W3nGOhTSASG/2TlIw0NUkVu0xCiaqf/7CfL0YbiWxBT
uv5hRViv+iXPlPL/fF3NJubEKLDACNROeRfMO5G6U3Q/dC87dVQuXWPAibuwtDJF
PD2HB6V6dxtbok5R9DtkyDWF9+4GrfkyawpxsNNIJ0qvDTGrkFw9nynwMhchJsJp
2teKoCmUNSYwL5FnSZZ6a25dENUp2EnRpKTA7xXhfbv+9L3jVZBQoIt1D+gLoupN
dKixLmANUF0+b23wYLqhGxZhgFIj1cqk4OnYRhlrqCLZSEPQnp9gHRqUiNLgl8kb
WGQH2+eBkkngOVXF7jU9qA+RPSGxj2cwpqGUXk99djn2XNwbux9qx7UtgLU5SIVt
OVZ9Ry/hTsWNGMDxebjk9he3UtZOCokL3z3XmFhxvZLSdDcVzUqLkuvJ8T5c/7yC
YC0JmR0S9jNG8/Ean2RPHpBMwqH98zztmprOsOMkkCrDrA/1wL1+tlnzf8G9Ow5g
boyVFd9TqLiCJF9ozqupyuk4qmq0FxsUnE4GXupRy4nr9/DF6gLc3va9tQNIEUFG
RFjqKwg4NHQeUosQ06sLA0S7mqNz/fm8XnTasmt/Ci58p/hr1JFdPYok2tUPFHPb
tuc94yXeB4RZ7jeGMB+BMnky8h3U2UFRmZKE+mCs7qcCT88EOs/2qXSoQFJ8PUH9
px8RJUkXsDnLBR9yUur5LoLfuyVJCcF1/Kr+uUGOhWl2P02ZE+5JesUjdkXyz+bX
cB0tviOg+0xmgpvUtHGebCTfxZmeNueptDXT4MUazzG+M25J34/I2zxE4+XTmnw9
1ohHyX507q24wimTP+eoMaxXSyWFsYoN6I32PioDQaMbdhoFhbA+3nHi5xx/dIV7
vhqtjKik5XX9fGbCHuAjgHhbcCUefgmAhB+m+zcIrSbEAM00hbaTNko/FF+QJGPE
yh+MxZVNjti6uPwpnD4drtiYybShn/WF7tMpsVbqezOUvDYmbK5QqOvQGFORx6lG
zNL0ck+hU4yNJwSvK30GpKgGta+5tKpP8uiegFY7nE+uOX5pQ/SDfY+iAYmhW7J+
yy7mmcdZgSasiIayipGoIIVP3m0uY2vt4ILWl01LgUgT8zygcPr/5Y6/FQV1O+ve
IhyjK24xZQYvtIFly9UGsSTaF07cmmnYQeFPc6wlS/N7Ie5ZKednEGt3/fRitIII
DzZaQFl/+I6BJ2ZOxSuy9avErgBtgrt/Ekp5fOkPqPBkXu0h2dIqgchgnIweUOdX
PuZJ1b5fkHHzf0d7XkEW7kpg26oTIOhq8T7kOh7/2HlinrK2ClG4nvqhhF9J0FbT
BqmKLznzMl0N650/XZvpzizfqGohEXXGP239lPE1armrNGxZdRbZ5DH4t13WUmgs
tzSbdMPomwhDctwrDBN06ms/9mTc643Hz8O0MV/tvwqVjbzAcuxISnKl+4tcKA76
j7KzibzcviCAhgUiIQO3DoJYGVnr17SDrw7uVPCP5vHCoZXaqauIoIQFWrScJMq4
0piYnFBG7L+ythIhBLxsul4X+0DLShqQkh5rV0krkOCVAcZnesTO6TYJlTo8HRT7
/q1oe9OmqJcocxEHZmy6i1k6XBtrLKbV5d0JGxHqtmZida98zfjCzGuvB7fzL0MS
yFNrwGT1Tx0g8ibwisgZ/63hCOHff+99ARFWldRjN0gftIwDiUSM3HffrFR5+vL+
mxbXYRaPWHUVgq5//dwBLnGbS5K3VRKKAGPbP4NAk2Btv5zYw7+FV/v9W020mqiR
sldvR9/+n75tzoIhdTPydnG5g7EdaL4MEo5Jb1Y4J0dq1VJlLiA1w9+DdN2zL/rC
mZRLMNKCELfxMoS3Jdvl1can3kmxCTI+hBYO56dEXJVi8FhSZvRHlbiAFjJjYcc3
wGch3BawhDMgYLA/BeIGKM4UEyvX840TKIw1LpNof0ZpEWMpwg/ZKHhzpxZMDqTj
Zc80dGNyJrXqR8kJ6LHNLtckJbVV/fJ2UzKRG4k+vbmdv2hcax66hCT7vByOgmV2
K5uH5ukypLoFiRqQi9HboA+9q7WY1BwCwbPBdP3bgCySuB2adjAjerDTirxXC7/u
HctPixN5s93H3VNnZxHVVarRrzJRvHde8HUOs79I8Iuube+t/gCFN67/1wQOuHYJ
tImZkMMv3bx3PGX69PgS6X19uk9GvMgMqx443YLXedF0Zm8UUrdOd8d+NkxOfnIZ
+1WkoBMyadKFlIvbceeiZcAv0sN8zQWYAoW6BpLFvzuPmTsB7m2k6KOly4/Mvc9k
BcmlxMXIw5Po0Xuwv+lRpB6MkRz5BQjPyoaA1urOQgoLUF1xRazCi/k46R3uEMMM
EOGDkBqtuTnJygibZzXFQ51kXGE/U3j1N3QW6UBoGudHOMUuXjcRobJYezkUK8ZN
xYEzoTs7CxKdNmKz1a3Ky1Jhiq/J/a6Os0/ROGlKAxD2SmpOcbSQRRT8dvEYPu4N
sIwkmbQkBl/Hn07+BND9l36izt2NjI+cmV5pWpBkgdAXq4kpF48hBwKmYDXbbDYf
Gj9k0b8heqJbo7DS5d4/QFfEaSi172pPAZeKY2uKFDTgFfPayVofuG6gWtWU2e4W
9CEa3W7BCELKEhEK7j+buaNhRCqhm1V/7Ik3Wr00LZDu5wEj+VCMtIN0AglTGefc
YljBOjfnTn5ABcfdIYVFmdsqWHZaSHXHvqgi8OVcPvYM1+oxlRFfe12zUFS8CTbI
BKhbWPgR2kLnqTEKXPUBdXiXP2A1I5Qu5tBnftdNOggy9OfNJF9gOpj96sY7BLa7
xDkmcq90eYN7Qoq42CbEUXsSUNY7pB8K0giijniNMALtyTPnKJTdE0NfFPNEcGOD
DUSEgp91cCXndVjwQo+pyZT0ZT151XygW4q2Od8E3fO/qGomhN1PyXN+/qUa42iR
Vg2WhgUvYQLJJnF+U1NxlJbvF1yc7Pgu7fJju7J5HaXaTXP/27rb6jRiyfsc+2P+
CR50ZqPkswkkuS656Z33djYD+XY4HlQWdpYW4KM9+XMctee/NbJYxwTx4E1q/Fq1
6DsYvLH3nyoLkgqiPeVg+dIRekA0IufU/KkH09FXVXXNOHLGIobfsoHHJKlPy2f3
VhRK0S7drVWJeO+W1A4ZXZES/iKwQt3D82Mx9ifYHCFcZScltQdh9D3XemRdY1Ea
z1WJf2uCNoKhLs9QirNUewN4xtZmJC172i9cD8jwmNnp/j/l4XcKJdYftYhWpN4d
t1sTUcmmXrqjEsi9TaanBUDy/HfT6IClVjuR3I9FfykI/VMyIn/+ywuB34QMQgof
VA1gr8GXMWMhxZmWmlnGe8rV+IYHe206F8SmKyl5HuZZypWXa2x6PoNWGXGB3lfg
f34YA8jiMI75RKknKBA+fO7LgqkN1qOAUP9JYQxQUbZ7bjVgll3RPkqmzV9Ubs7+
686d3kVUMMvZnxCRqDwvFRLOlagwfB5MD2hyncFtBqKTdFhNyy15cRoCYna/fR4v
40GvOuqoASk88I5LW/b6DwoubanZge8np2ybdpzsjmIydSwbHUomQp/Uw/CPHZAo
SazDU82EQASEOIF9HxOj6AHut+8ZtZeYH7KREUskWZGzgWieKl4MphHmlrtZm9QO
R93ceR6y0QBpuaobki997Sop7qGynQo9bKpmAjw6v4TCqEdnaSbiowKvynupEems
KQ8Tn6g+d+U3e7wVnxHJI4RdNS0KazGerU9yMGSs1fUbdvr7ifkHHrO97/vo5h+N
h1dlE7c5yeK+751F68huSDrnK5ZoZbgaXOhjWNLnNKE=
`pragma protect end_protected

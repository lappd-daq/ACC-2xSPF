// Copyright (C) 2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std
// ALTERA_TIMESTAMP:Thu Sep 13 06:32:38 PDT 2018
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
GrXC7znaBWTa+n3DRQRMY7kCyw0jfAQeJGEBRYX5gCnFKU0wf4FB46dtqGMWAm4X
JA7xA6MXfOT9NsAUbAs1H+jUTIBt3pj7e8O7b2IbiHf2yVlNovGYZvfjjvdqss62
ERQECJdNAX4pMVBmnWQltWwMh5ol7VbHvOf9zU/J61M=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 15680)
H/4VNVRwyOjzw+RKKy0mzrEaqGZLtZkq0Fw2zzaxcnq6aH9nu7IbXEj2NkM2Zh/w
KttrZUFEMo6H2WUSohqDD5G+/fIyAZCcd63vkNM+bnPuwp+BZljL+maIB6RZMDdd
PArpouQ2M6uRkV+skjZ+fWSrsYLNpWd1WCEpcr+US+bwQcj0/oeywkCKY5wdFGuF
ySepayISfchJSjJAJK4rU5LZvvJMEHBb/efPLSxiW3ELA20Hxn2Z933f1EBTqL6I
YXxDbKPZuai5NpoN85CSsVeDqh6rx0Hohal/7ri8rOCalTHdMecRxrS0hxoxXM7b
ubaiYmaKKyq5R3jHvFKQpBudrzd1DkzXhATas7BO1/MniUv0Myhnj4AqaAcH7mLU
GpEZg+HXmd+QNE4aFzuN7JJVeB534CO2SgP8B3MwFiRfEjHNL7XQ08X1n20dkks4
yu3qyn9nyhTNudItt2PG1X4pA9uGbB1YT11fVBV2OnDs7WbX8p13DOM9CZj5Sbgv
qRHjVwYZAoBy4PCdfYF77LxdQ7DSFEugLBTIsKMlPYU5bIbhoNyGqGvG6DvXbuAb
+s+AUfYJVEBhdw/5sjV/M5/IZ4dHRh5aGQT7lnIUEeEVb4FJkl1ga6JOjcK6C0aH
kqu486qvDJVDkZ1UvmY4vVGaRq4EtkptNIwjF4ni6326+XWZjxz3ZyUlA0jyYjl8
kgXqT+qQiocvfljpE/0EBIc9+d3C4Ndu5XO67J9+/5RywabmauhtDDy3eOfJk02y
MtxpCXChRY35JfJmECDW1VtMIGl2o3UyrY7J0+RkwoVm9aK/cy3UW80VUlSO+Oio
iJsC/5fBK6HcZ/Kg4/uI23A3zJArQzT4jN29q8DiLnLTnnZm0J+aqApG8deixqOj
OcdT1DDqBmco3mjw2oujpNrj4ZrWXYu0FGgUXQqGjHWIovK27vArdEgvsZ63UeC4
3zt7V66pSnaTpmNepeXkmxkcWpKaZ8lk5EhDlqfNr3BkhrCgMFXKyW7eByt3Im08
sFQ3X9oAhLo6kjK6ahsugLQskdGhdxpv5qsK0zTv57T9SyZIbY3EEKJjui2aUq4y
42u5xrYZ86Sy/mC6IcfIk5G7gcQteFjkR0qGhcstvXRauAWd+050MhUQL8up6/LH
scqdK8fULhkA+TGRdzakfFzBE5A0EX1FzMwIl2punRRayKXQjL6Y6USTUPq0kA0s
ooZiSmX+j/ZItDgZc3dikJPBlxK/XBrQQ4yxBUPDXsnwFaIvZRpdnuMbgmBJxds1
wBKaLOmfky6Gz0iNbMBVdBoqRU7XIVAIaJksJBusPP9xg2pKbajr45ZrigbLkAQC
5VIBmXEkh0yLjmNPVPoHd7R7HgA0+vjxIEtpb2GoO5cXmpwg95pRVcuPG6fyJTzt
Vd+8HyuZZ1I4khipCc308Xygd8tBArMaPdABM8qKYDDLpgg5pRESdNcKMzbmKbiK
a6ivy8inlnpxqCl82JPVPx8MKe7VpkGcaYgjZRDvsYwSgy5fmEQ+6olhy4igKirl
96KEQvD7/LOwX62GWrJ441MpkNx8M7Q9riiQt/QyWxkxAMgxoIWE7EPlQ70R+Pgp
3gVRgTGIN1P7AbC49jaEaWI7QCpCgEFgF4nVeOdcu0e0flfdKIUONq0o3Jxkb3Jt
5DKc5KSVlsclzC1YyAIzzpklXqQvTKC8lygWH9PAW85MilaKKrgfMkPh2yyCIIMq
pozeBfVp7uXXbo73IFK1eadfHjGaGMf3oj75XZSb6Nh4o0u75AF6TSN4IN7HZngx
aSOv7UVFOH5rIw5v2BlAWEgsp8oQJ2jyjg6+yJZ5h5zst/F9xkZnWzVQe+sEiblT
knqD8rE3tMO/DxZvDBj8uJIpwbL9AkWaOTI1bs3gqHDR9ek7FZQ72rgOXplqlzCz
ip3ZlS3o2aCyweqv8Xg/4VI6GWC8Yi1OmBSlnJpWoRGSUtgE6P/yhVtvlY5rsaRF
zuzHH7+Ccfztz53LWf5+8S5VnbQ7m/v5te99GjbWMmRbOOE9dsVXNR9AD23NfHF0
UNXo6xEOsxWw86hB+Oi+h70ThHNEupwNuohsbsb9g0GGhkcgzAaSPKjQZhbok2xq
PaPCXZb8DUJ6isEggmZuLIjZGi9yvunBN5uo7Ij6bN6P7GamzEgGjsPmyykFvRqS
QeRFqS2w3pwlIhuh/IfPj5NSRAd1DfvSWtaI0r8tuwgKL/OzDt/j3J36O+Uni+Mm
1EdLpRwU/gSROPAB39JjMlRjTX1rtPxMIf/ateRgPndpFXiVijvsfAtlvyOlrFV1
eR5aPd4ybeiMtbAeOh6M6iC0R9CojlfVNL7y+buubenP9CLKCbIl+Yw4xRctR3eb
NfubHgdTbVIb1HtgIX5dplTg8qt8JH6GivjD42QNL8IS2mA5UtRMV3NlIO+NT4MS
MgRwgKzqcCXgzV67p0xOxyqNNrROrovCs+gVDx3WphjqBtpb+KxttS3exq0jL6xM
x+6fJpJM4zkvroNyXZ8REmxbWh3y3/g4c4uq7SgZr9d96tBJfj67cb5m5EQHnfkF
80yys93/IOKcWuiNYfPXmIdZWpHZlCogdEHz51volmxf1YlBWP7zut2/37+k/BfZ
vIYAQBgAFvVH2AqmJGzRBiLUicRmCK9bUFuiN9k7bFXTEVqhEQic3xfuVYcKRn40
X5GP40652VCxwn8sy5WjNvWCDMjso6D+uB+zw9Jusv3/RRqo5AVUY7UAf36xsHxK
j/1Hz4FtZt79uvVvF4abHP+1yel6S7Y5IGYG9b87q8z8lOnTBpSzqLLDoCJ8QQAQ
Vm1Fwq31j7QUAioUxN9AlJBKi2QKgELQyFsNjIITkjixNY/yOTUNdKU0FuKounkD
nguq13gZSi96rrum6vM3tOaf2tpRTUpN9bWQOfGEzwoRrm3qGi1vj9xqpYXxS/EM
Rcz9WPUdvZhcSZ+pjtScaW+9mFz6WA3FUq2Dzh9DzViaztOksWcJ1+U6Fimhbraq
y4BkH2Zsz9fMQzsbPuGPXkXpaWoG817ijTJLw2iL38uNEuWnwKHLV5+C0lKvg/mh
TpugVnYoM8+ffbJ3tE+SjCyJK36BW2hvzkWzgQkUk/7ZKBbyHpuE8UAPyrCAQqGP
XijF+MBMpLCIZKqCmv8UkZjfYYifNeyyr/UBZhmvux6XrDNdEj8+75NTLSVtpXt9
j3F7hp9OxyLX5ms475ol7Tq4al43wGMbN4rg4wwjsYwzXZtaNGr748TKo8NKvpND
VjbzRVdaVy7YAIWqzBITQ6Z9fpgz9kcMIM98q3YK3nuagCPPjlWSroJD2tRjw76T
5hkAGmRzzEGk5GJIcvtUidXPlBeNlyW6MV339MUCaVrhTmKQdpP7FZbW/kZ9nohp
0ur9NZEHGttEYkyf01yNCDc0Xe9RWWGj01L4NDc1roFT9vO+uBCHM5oT0QRVaC/C
4cKRgi7Ylxz8rVxVCMCPkil2S7cWVTbvTSAreZHZDVjUS39G68EQr0pZtlsfof7p
aUlBfZYNBsVF1lSaGqkyMMteFJL9y9/T2QAE6EXi8BX+zaG4RC7k7gOg3Zp+cLYZ
2tM/gYqowIptbV1vTuPV0U1GJOds/XCbpLoPY1Uw9eGAXeRdGFNUQbHJ6KhRkIhz
scefr3QSpJGE9JX6PCPC3e37ReKtU/1NFDD2CGPRXDgZFkazypcsffzfoEw2wMqp
mjqKZGET0Ub9mWNjFj8S44vywORKSyABIw8oODBypGqOQaHt2YVgtaUo+DtI4EQI
7pfYiFnCMYL783DysckNB5+7kF1s3OyOY51oYM55Egcc6+EtGMYwK+/60I7MPdf3
Qnl65jDDsrK4AYQFZDDSLJKmlV9FZrejdQe9VA9OElu1RWnNGUZCBkKbHsGOlm2V
WDIic+qGlAEDuHJHrwQthlYlm4AadA8swBF2maKGqzbVhe/wFKoNwXtD+KNDpNw0
045rUS9tbBntn9XeIV4oHuyOJRhsnzeztbWJiYyPAP6TBHZMgVA5pN6SWA+fE+dM
58GgFlqj24ERt+Z3kLlVbPmXTMNonhxc2cgKTAyhF6wBJ0orEypmDaw/M3qq+fI/
RsNpJDikbALPI9ivrPM36lRgzkieGZXDb4YkKBEjEpg9RZa+F8QOFE0BaySooYVL
n39SXfMTwPXGTq2u2bWXdc3LCmFgEK/c768Vuz8kCB63ZDNYA+H2Zkj4xP+AqEPZ
0K/cwqNlU/AHmUzl6cSw2mdDlsW5JSYH2GA0elsAIj6fRT4DJMSgdPWyS1blLuMb
MQt1WSnxEA8KFTG3smbiA/W/PZowmeETLoPJvhmfurEPFVrh/9acI1ljeLibn20g
qUKcNT2nt+5uuQb5rTDlnPnozjSHuiZ5G1fUYR4HA3keegbdKr7pxeLotTHZIies
ScaGIDK/80g9gLRl5/SW4V/joQBGPZ9D2MN90g/gPyDdnPH+UmU0+8ijS1MFiCWm
yhcz4+76qRP8FssRUJAuidhTAwWvRwxHX8tD1vpDjZoG50Q1+C7Rdj4J8pJvNNiD
mT/2BFBZqbt3Ce8sk1ASAtTGe0m0cZh8wotwP7d5gQL1sFqAxwfs/IJeVlbwYQGh
ShEkv3snCOxYgSzDq3xKm4zQ1Doz622I5BqKNBfnnyye2lMo13hfbNru15H3QiJJ
kMlz9edOi6tSkqPlZs0x/7dxC1hkg/lRpMMRHDpbHrOW3AKXDpW+PUMNWtrzbXzu
7LQ13XeJ1LlqThIEQ4hUd09NZg3PupI382SHpFkZ3NM+lI5MZLiNUZ+Yb7O/bxsL
QYwhcNmY6mYmKNDYx3p7yJKNd8YR3VAiXas8soNN9q/yAqUZBlEKAAB0yK0OeBou
Rqu26iN0xvS8U7O0Q0mLW0Rbn73+G2wrowDNbPa0zQBZfVS3l8WMzOywJQcQVb8H
95xEPWjzNTKzlngGQRbjv/gmPPkdJa2eLodn2jthPuW9hYxJ2PedL1H5zUl5EQ76
1o9kwG9VU1LvzT9mJrIFA8UlU6ztdtjHInsu+3yqCc24CGP2Swul7M2kDDqBdJ/s
2xZAbjTpij8eaUTSP86OtjA/qsDuKCQdRzyErQMq6G6OBqN4zU1x26JKQ9XmcpE1
DS5ZyKacLQB+3I8FRaiwZ6yrzEAdbFI2p0qoqnZbz7DW7snmeisP6sG644P+Tt/u
SESiKuwxzXiUMs04IB6eHc0hFG4lhj/ZPG3+ojwJjLU6CE7iLP126NwLfescdHTm
cIKECuMBEoQFP5leIW3CoRVeuBQV7MpwKT/k7t9aYQ0UU8evp/TUakGckk+/WgRR
/QXJcGVlT0JM0/shwMIkWb3rVnRXi4jbQ9S75ZMuU/gh9a2f3TpR8eUGwE3FnqUY
cnAnSSBLYjoU2LnWSxH04/g0085uzK32FknzC1ALnIzfra8h0NSH+w3CoDJ9nup+
vr2zEDDWHQIyL15nnG51yqePzgcjhXfRvx5tAajDCNdg5XZqxzjje6gTcSjID19z
HBB9sS5vh1U/2jT711WFpvNpU1/MBbz01ofl3tJ/FFhThU8RFmFkyNFMh1VBlE4D
PhARqj+ZkCG4ciQObVDwHICbACkZj9X5ruAQKJeVGMArIJwCRKNljpSdNmknvB5c
paPibuOdAkpRK3ncl8jzhsry4tzDZV94sxOJesc618nefFhJVFvyCK04T8vEXC9C
6d5BiLrEpgjt33uuqPVrkEahNWLzowrA51OJcF0KtEBw0t+By0dQyhIe0TZucmLe
/SAPFZdY63lo44ZhV8XcfPOrjyCKmjFWMt+jzPi/oxZrl+7BRekz1umN8IRzxWiT
pqEaP0S0dYri8mbhWHttKStVZLJh7LrY2kpRes3il0L1il9CfZWYvk61M/yPRKWE
MsFG3Q2gcYnsXQ25kCs8ctnGOQ4l1U36nAOFowmwjjAE31qt7iBq0vE5iQY/COWL
UlDrb+SJHJTj0wa99zwVemcewIuCxPLBxPKcVbd786IYkiebGQ8yASC9oBTnYYeX
7yBLBU5GTGXozl98MB6fdryWUmqzunhgSzLlyqk1GD4RGAnl5OQiUHhJIUSzf//Z
4mBtkSnX25C58x7VlslhltebOw8Q8z87eIbBWSJMF+7G2lGesqxzzGYH9uiCRsgD
9D+Z7cadZHPgPHxXb4AG1+DkCmznj+4mG2eaQOW2XY9HyBHXaVnM4Z8lbJeUgBHS
Io1FLlw9VCNquyw/b1gskCREgLJuoM2PBZgPMfSI1/z65NPDnrXqKX1qcUD6zoTF
YEOsfmW4VR+dPmPA1DPFKPeYzVyvFfxhVDE0mVc4LfgKEuqwYz9+ftCP+5xpO4wH
CLLnHdkQCNNoiZlW/tSGBDeziJshP+8wV0anDN9nyVMd2PGIz6mo7gIrb+lMBpr5
UsOa0h6s/eJ18QlTtgZ6V1oVaHKjv15QwFHgc4o8BY67AJ0H1DgbpelT3/atx1w4
Ywv/jl2HxkSaR10NAoCPKhs/rAPH9kZXDjBCAFomrN60u+Guwg9YHyQvd21pEQ+K
jNaGYJDkyfeHacmjCCs/7wZ0D0FjoHcmfpu4rFTWs7dtMFVXaVYaPnqp7ufxsMKT
W7XkkY9Nt2c7S7NB2qDBd9QnU0Zv1/1v/rIempeDXWKG60GM9xiutHrknZUdj4PR
IDEaVot/UIFsrHn7PZC27klbxLbTCyRXjRwPTmFjI/EtZbj+a4Ai9+HWPEXv4jM6
03lqXn3d+uIu+TaoST+Xmt/uiFWsqlkETyplGMk1zbdpXUbitKtzuXSGxbUeR5OT
TT936+3nuYY41Wf9NuV3rIN5q5AJDPf3FGGfoolmN8xYUcOGezqwvDre359TuEFb
M+RSVnctCpY9ZmnUxBpezgZ4y2dBmmwuguGCMaPboKE/t+QxZVIQ8bTRoPtzuGA4
TKzV14jQebwge3NqPnFl6bXTnRAIidCE7QbGgS86LjKLzHM8iA8CE5JI8HYDATN5
7V0IfK/QYGFbiWiYco3HHSTQVRCa2hRcJwL6acEOiluCg8Lrpqxnb/Mee24iH8/R
sUCl5Z+LXLtq++g7SyeD03Pc5gL7zvCzuHR2jWO3x7l3dlWyNnh85If9VnINDuUe
V8fDWDiHopYB+ZdynIFJa/0q2z5Un9Ph8IlTwZn7rsu5mFxvaVr2pr0MopbQXXML
4pg7qpB3QZKZge4TTY/d3xM9Ddd+x4cNaP44QrS9ie6hCxpVoLlZOVK3OwWjQfbc
YpuQtzQCpIaUWIOcRZhjy/OcHlGGuKe18zFGsQdvYmPBt5+WctucqhowvsD1xeTY
b+2fSr6/lmGOp1397wxKWgr8/SvpT1Is2G/fBfnORrJBJi1ALP7TD75mGHMogFzY
EcMeX6MJD0NO5fiUmoo6bvZnk3dwBaHNa6czhZ3J3VeQA0rgzC+Pgl5cDoNDeRiK
LqoR3tTPwX6ZVtjdq9RRXIY1JNOC6ED3uiRDEIb9uG+RG2dF4i/GHGdG1U/ZrGU2
xmoQvTXKAXvR7yhVKgQ0F5/tcXfCIlpX5LwvMNxXYomFT3grgphpXFT/V91zmIlO
sqQx8BXISIl59RpsL830OP53kb9ea3nEpYlEZV5GKSnFVOpV2rEqFy00Do+WmZnv
obisYLVnUhonmYVCOxCKqeaF7aSBtB60XRhxraJY4EjUuSLGM4FqW0LmlpGPj9M0
gw1ZLIVZHd8XgMyFU386l8SCBhispDEIaNlQPdUTKKZzSf0/hNSReNyARqbmn3ah
yaDzF9qDlYrRzeqZapygTtUOBdDOIreJw1f8a24dky2xJSu5cS8RuryY3AgeOEac
D0lNhkDIihvHJj1rX8wh6iA2aNQtntoG3f/L64h2TyzDebSUh/tS7P91AhCayYaD
x3/YdIjz/V93yI+plwqzdg8TcW0PrkW/1555DKPf7BTk6He9H7iRXf+IX7W4JcbQ
VK8TsNAU/Eoze5RIXQESvoE8skMhS6qgLna1FHa93faVIK9U++flRAuw4TxFutX6
nh+AR/1n0wHOWHo/AClCZQkyk6bW41GDtvipuudu4uHyW9Bo9vCSOmPVc0sWYr8O
HBEEXuwAMchlhjuMgcG3NxpxCAzF0erePLES1rtxWSMB8kqkyvd+vk1JSTMzdJzA
PJ7CchwU2FbT5sOXQ4xaGB5v6+HLmz6xXZ6NvZDArpvYkCzs32E75/rzU9UoKO+D
XlVrkXA4adIGg8jgPh4bHSAVNPPTRFCZIuF22QwU5z6rp1GCqwQ7Ir2LdGK/WG0I
5Chu83Noqr1kurA2p7T7zjvRWckqxO20kFtHLRcbjRdrZoGQdCXvVBmbtAiqAx94
3RPpWhD/goZF2YMB1EAa6pPdG3MsFsLHLzkqUsMDrqC+AeD9yfXFNc9hBjyQ1K8y
WS4jkIwo32iM30t6gwtDkEHPzszKsxH2q7QDBYYrgnqf2McbrbiKYIj5jrIlaq3W
bjoU9jilBGkTdHc3QzfCuQI7Ji9WK7yEwTji8vCb2bf02JRIpqb63ASbLI7av7Zz
M0Wz6h48E1avvVyYNSManGeqPu2fe/AoLWKyoHD7QyBufe6XwsorXtVzQJMn9668
ISG1DsSrHeGSr8Lb+koZKxRuCFQry83cDaJXSjT7mI4ueoCh66JYj5GNP4Jza5GK
LeOFEk0F45URH4rdHj/ML6VTukyjAYpRv2He+NLoQZTrL2emwL/F0Cu/H4xV3Rsa
yEJBoDB8tYhpxVigzxSU0Qw1hlVV6ITWnw1gb0R893fWkBrkumjF2NCO1+aaaeVo
UMIe81MjgwAkZfQmDLuvId+t45bP43jMqxeVNBPACP1GgamHDKiBibiVDpsNOdqA
mSkAzG/JCepYD3yXef5dNtcLRKT6PCcu7/5iHWbpLf10vSveAIRn4nJ1pU/ldx79
ZpFskjKfX8iv2kteJ2oRHDlej47wsbwA4z2WPwbR3EHJ9Ey+QnJ+NppALGPITRfa
CDAOSgAC1T5JKKSzlqVHhJkTNXgMr6kYYdw3pw8VGFbxe13HMmnVopV1qzHV/faE
umm9LwfUg69k75KmsKTfV8dFt3Kf9n6t7vvFidVz6V/9ct0yL9fWxNbeuXJI2aRz
0AtgEC19xV60nCPpt8R9liYmyfQkqaTWqytbkWTOcSrMKxQFaYjrSiBJ5S7RkMWV
p147zQOZcdoD/2WeUQegUPSUFfCIywDpvPp0iG9kOZkPXJNUWxPPsoPVpzxFY6Ns
jsLvMmpjSVESVHEYSrMy1/4jwVS1U/pxdmk8jNEbE/vhDz7Dgz/iv0qnPdYqy0EQ
6hNTRwmhst9+7QnEv4+JGuNzs4tq381EXvdFMtKxYnQ0YKU1Je50W/Rao6ieuOZJ
ceCxXzLEzX5ZORwrzGwjLbIvy8JeqW18fVZlPbMNAXG6Q4BX9lkwUtQglLbQwdM2
zyJcdejnErFvJIbWvp2dyYxuMuWo10hhK2oD54G59pQQg3OkMp2sQvzPu4VG39BB
bP57QwPQGwFecngGOsoL79yayBb4qyIjsBdW/iTCgqG1nrwOxD7hm+HoI79WLRZN
la0to/HSEy2XLF14EsYjXb9LVR1dlakbEH8Adyrpbkz9OseqEqR5mY6T9auAGXLh
+HLwpbFHnPqGxX/Aw/gZ2W5fTo7nlGG30g0OqrqZ8li6Ixjx3lK/3k6O4b9IM2Uk
Mu6soWGd30xgfqg+gHKGp3xQLJKMYGFtBI7TOAUgK+UEaYu6DMJbJDR0iPwUEI0V
IxyWyytgKk54TdTYBxfzlyuH0nBa16gumnUvUm4KedyAnBkg/YQZbFwzoU5TRL3J
nCdLYpkbv7qP7VWK183jWKaXb8lfmdf24SItD82q49pvrEHosvQFzP+fdrEidX4t
FM9K6Hu2n3/f/FWcfzYUd2wQveL3u8tQayuaWgf63t6AdqBm4ui/DAP0+m2b0zgt
2rhWUfo7+xpyKcU/NRr/VbfTsmh5BoP6FAcmAKkR5jyxiR7wl3HTnDIE8DoOkfbV
dnwUP6hVfegVCvxQjMxFY0xNrr9QAjSRsAtFs4m82PyydrpTbvT7KNhybp2zahxz
4vt/aOFk6WWrE+Z13YrWDzuw5I4u+YLkdlpDHWVpWm9ulov0R0WeLdXossZozWWs
e5Fi5Ejghpgh/SMSv+6XHQxcSHVAMIrqaVWTDvsrZue6UYnCALHbpgPLw2svAx6o
jNgWWxscCT4eQopArvMm/PC4t8sfrHC2GqqGOWHAPhI+1DLLMtdOh8ufPOU/EOOq
vSBDh0mcyhJ14szRSwLD/Ka+DUXMTmfnQk9PaCEkCK79dPXevbnWFel1Sdl1l7j3
F9TiaktYVGF54qHEWFfXeAC+7w/Y5ca0KlzfZ6mASh++BaKSeQ7Iw2jr1VGoz6Nt
XO2EA1rpxksz0LTq5ijPUx+Qfbc3k04U7pO2DC73NC8o6OakYvptc4zTvZMqaAzG
n7coVh6X/lm6bOzj8IXxZH/m0bUKxyceKJG/IIU1arG+M6LzOjeUfTdIjUcIgAA9
+oMnnLMfxK/dADqY930qtNfPyfwAjjIGSHRTLhEy/YmuJpGV0O1gnLsP4mQISxqP
1QTSU1Dp0uLB8L6/ViL3ozAr7oesZof+OjW9q7u5TNufb2xFi/jW2wjzTvDMdBbp
CT2/iK8UFVI+In8riYrrPbKAKB244UU9+eHO5V7EugI4bRRQjS6txTl2X/x6G/EB
zVUCw5v40zEewCa8lDlOBC5phbTVhkLbVAki0yC2xClhQCx4r97TPEWSCHZkNZNJ
mCh8jy1sivtTf9b3YJN5k1pps7yJ3Gs0IEwYKioA+4u+sVL+3E+9kl41vOi1Kuyy
3BOSgaE2Jq/5QYmuofKADwak4wBv8AnR6CCl+ZumKb9Wwhipe7EWujVrKxHWe/o/
CnXKbZ0KICnhSI9MJMdLrC0VpRR0pHtr55Ve/45ZYTTgyWTxxo/pfwD7+VQaYeln
Zw0/Vm4lttXeJa07lz4JwU//y1VFNqwV5L4tf6EB7d5j6xPvIwrSXzJtOu606v5K
EEEjWmyGc8W6MvqZEKNc6THqHfaQ00pcjMBNKYJFelFLgfB+QnactmhbpHdgzB3P
bjF5t5azM9Bxv3wT29UjEtAhshDVJ1YhT9uLrqJZ+HP2yLN45Ou5m6/gFXutGlAs
nluDpFW4qZ08oDrQGYPU8kVnIREHD9til5QAusNJya+X3yPQ/+d0MVlJFIy2aDDl
2MkTD0S7yQvrIMpnpeHloc6uzjIhriv0e6qSPV9FiKsqDOq+N7Jf6Vm3OEhVbAds
ekjjbgM2UdpeKIy+jr4uKaBp5q92bGJFFYdtXKVAW2ruy5sU4OBrRtm4ExNTNacx
TpIMHxV498iDxcscunErvc5VgDYh2z/8h0z7Ozox5uyhlerPpAXTO9tuDMKHIp8q
PjVyMMWRNlU9+bruwEXEHoOHSYR3cvvKaq34OOAdPuw4yVrLWdUQ94jzXjE+RwoA
e0P2PbvTX6jgXjaN3bQxl7cWH+t/izOGJSDA3GRpn8XF6dp/9tqW4EFj5R4Al9Jm
zqB2nKj3p85pPCW4DnCbZMWFvr27OPA99Nkjb2PQsEDc2cVcGWRPqi76aDT+lmFP
jmEe2sy6gVsMbLgcOZ/EHdj7gy+jjj2/szwYNWxq6iE29dFe6YbN55nv2kMg77p/
8GK7oM5LxpB6W3Q6fyu17aPE29vQ3bBIUIWVYlrZ6J4NwC/+mIOxLCxrtpn2Esma
7hwJ2nhUiFPMS5JiXPh3pJntmaxIRYktLG+cwfu1ztnA9Y1a9721njbdEB59vz1H
5UqNVdRVvDg8y+jnld+4+w/OrCwU7ZmTef0od30J5z32HuNe27k9K71UWOOJTmRf
pqsH5PuDayC3gETK4hKXBIo3e5HcOjGsE4zTu4Nu+E6E36KSgwOzsx7RiGqVMWNC
uK6um55LJjfdyJwI6YF/GxGWtUxLw908kvbl45tQhJcNp6GmB7Pp2Acy8BXqDBeZ
8EjcM5e+qNjW1S2w9yP8Lax6Hys6Ess+1hwmyBrHOHy1WrBz12XbY03u3lElJB6g
2myzL3U/TtEqp+gP5VlfVaHooyTNTW3yXE4Qfp1dMWJYaQrNmrRxLZmpjmezclcd
qNQGP4SpHVfu/g7zCMGNLQXOPYjLKenZbSC11MOwWg7wz3XQSBrthXioZ/e/2fE9
LU3hx+6intCI2jFec8JU2DzTHjVq2yphqIgp4JcsRRp2sHT/qXGEhGv/NJNWzxfu
ORS/N+NZdoG8xjAWGrbPh6SwbPQFyW0OmpMogvV6DlfqJ4rQ7CCfuRbn/V4r4ove
yc8XcpV/LRvb/09W+0Gch7OBD5HcJxtrO+XqQoK7Z6cbAxzUPQEdJ59Na+5svk73
86kt/BS//rMQ/DAydKu1QNOxilGgAiPe9+u2JeOOxINmrA/TwxkHwrTKD5HuOo91
N+GhuRLKNMo5a22AKDlANoeR/oaVNTZYTxMTL/50KS/M1hRTBktcj8jHuz8jqy+F
nDckGxuffgULgKwHuini1cIchBLGW3/6EOKOIa6pEPIJfY7lSy+RMqG+y7X4oRDI
JGRAvLQqzAwzsyz8FdkBmfzxdHBNIVpa37dIUKIO9yonyvSavRYmn6voPU+zUGmc
kYkiiYWvtUJ0VsI4G4cEMZIEvx+TOF1GOyumafb7LVrDL+yh3A4LfEgRLY+aJlfZ
dQNo/YP99YMrq03ONOURi4xL56Qj9RY/VoS76Yq60lTS/izUnxMfUXZRCjYNJsoo
1r9SSDYFI36S05Gf6jW4GAOKq0Rkfpjz2lDpFhaHUkkv2WUi7wa7O42cjcVUtlwc
o8t1Ewcc7DHYYYtebyG+wF8gnjqJdEF/5WV5D7s/VWvd1BSBmZNp5LG/RMxw/24n
L0HJUzolUN2FSg1Q6vBuvPz2mUHpampdirRCJ4ZE0b6bmvkvfLOreaYUb3J3uoVa
mBeZHnbM1BSE7B7/MqhQ5WiP12FVvDFH4xuJlGNLwmLKXg2NHF+4HjtYkxLDZTq2
C6PPQqu1G3tVf9rMk75TMP5TpL1BEzgZRE4pBXd0b8JMoI+Mr+tH+j/e9aNhSiT/
dTFr0t9LDAR9+IM3whyiw4adCzAwwNXWjvaYy9oG9VPAf4oMIYmwn4QMwkJ+Cmys
ydOSrJ+485ZOfn5Do+4MT1pN/5VKORCMx4O+HazWsrKnMuodNxoREZu0wQZLtui6
6qJD/+4sbuAWxHVrGO8LIaXDaZf4RtrXHTqSFjd+CHV9YAQynx72htKaMl2stskM
eXKiBkThSrUcPCGlXwGwaF8l08rbebxhb0Onc1eXhdRcmcXaBT6v7T9djt27FuLX
OUVNd4Uah4H9YG4Hdv8xlY0I22CX/fqewiXcvHvchkeDB1ArKvu7DfcjR9mB8dlu
AjUjxBv0kpOcdiYbyPwlub6QPryojn+G0yA6G5BzLeJVlTNDJFVJ6YL6Zz2Sx0eB
M3go1hNV1B0i5KTpoHLM16LM6cchk8HloUgeXnPWvjsF/qpZRHrXl906ioKcMI7E
FDnLTOcyG/rZHwFojAb80/VREy84HJRAdZ+K6u4vU7OOckJjgc4ZoLWZoxaq8AZ2
2c9jUNFi/uvY1tswJ3nwubJPoNZzYefIlbt5obBLPIhcGiyoP6BDy6zH24mJ7nW/
GM1rl49rXDSlbz2sM2fKY52Ii1GQk67QhW72skTm7RetNCIlSStwgBUzWzuihPLk
EKuqdvirE840ddseq/yqBVlxyS2W5uffOIpdOJ9I42N7eSFupy3VtpG8ttf4xHrv
JHOC8TplR4adVjBrxoH5JIknKlhLln8M5Yd/fhxZZYrP+gZdb0soRemwGCIoO5Ps
fpWSUBnT/L/EiSDlBxehzgmHsTmSP2A3b/W+vLEoj6H0LffDu2WNYs+MF7T0t2/8
vGTtGmwk+0hYwmnDpeEXijJLBqXrsTfKC41RbtK4/Jsd/gk1OqWil96+s4i2rkNE
fVIJ+bJl9BV1D1a+zMOC9Oh+FbgCKy7h2r0F6DLgkefrHtZrJVmh4wpHEBrEzpqo
Kk9vvSdvARlZSKu21B5TJqaaAO2JhRKm7Y2cJBiUKZVxLYX8Esb6ng4VZD+wcfN/
BvAJQ77i5Uxn0R2yCKgktTuxyOFzHU67kzKVGCNFk0BUjvfoOhiMHsrCED7iETrT
97PFwaogBQe0WiwR31Zw+EKkcoO+VvAVJ5GK639sDp6mCmHfw+BVCKGp8+fsTCRk
T+AjgqUa6dxn+M+3FblsmysddqZjKqf7cDtOTIKkFiKzItpnmcXgy3lx7v/OsiK3
mCWDo7rM8cGXdrVpDKkty57MuhHdlogLJgBhTquUgmMKUF/Tr53wO9O3KYb9cSYZ
Ub0UzHquzoiFt2Mqf5ku4rJU+6uO6Y421wwWFUsZWe1iTVc+SlqC/BZShGA8lPzD
OED7kUOxNzqUxnGVjJ6TPaDw1vqyPYP/WHk26Nlqn++/baM9zHV1Jed+g22H0pzX
+cOvvG5gPaEYQGWnXRrN8qvWpB20dR6crjz54MWgLQVkdaWBrAtQVUnUEsIHr5+h
tUJj54gzb152mwJWBEf0Iq+StwFuwPxxoD+Y98gwDuWfKltIxTDYvmctg4uxZP8T
7PBsrurMus/ytyrhoGqJ47xmJ/MeqG5nNsL6Q95SD9Cqw4i7xqA0wP3I3HQtcWCf
W+Si5vpUjVUbZ+yeOGQ3HlyZykVIGponXhknbHPg1WDL82Er92UHfXyTe+IiWDLH
Jf0paUoRv+gZw6p6pRe2BlqixlzSdVDxZrfpV7y191T2z04KV5rohu6dGOikxlQ9
KKXCD6GKREgStjnxVtP5nw7zOevA2LKc/x2bc0UO3JOuRfq9Tajj4lHgEYCraTK7
w27LHUUaBV3MQFZRH/jQqIsbxf/5S7X258l/MmCMEp0h9QJ69SIDQDnS5535kOtw
c6bMkNgH5j+Vfkd3d2HNGSwVE/dLJFizjN+h5uaAV9LOdReqe5li6MU5JUU3B5us
pe4w8xkfaylgLbLFBGbSHctMQNTt61sz7iVbuJ+dhFGe0oUifHNYqmfhILXJLt4B
gNhDOhTomRZSduPpq9vWbweJphQHBXAK1a4ldVEUqu4jpQcgsWs6lIQN0NsQ207f
FoO6mfZ+kj+bdbBwHGRdPj1YY0HNleKkWmuWFs04+OdiErQqc4UkbVhOqcj1g8iJ
jb6Uu689k98c6zQkzJEmZvvgzYf2VveRulMPz3CK/xol4TbFvm6H6E0K71g4eGE4
eXt3cCVOnK1W3vk02MxOFUqpvghwNmeoFA6SKp/eAomdSQGLz1iOjPWr6P28mBcC
8hh3clSA0djCw7yjIMn0g0VjnYNnA6YCZWc+YdjPe0xdIHmtOWz7tbL54cRPVRJn
SVI+eBK/vkwMvy1kQPiLkaqq7LlPk5YdLcgJHLXuUoTONPoGnW6GSgR2XERHHRtB
c6yC3s79GMyKhabkVCX+f8NoogQw90WG8Fmkx3oq2PwIkzmmPtt3yhnXHgUMCqfo
fNgWGMSeQC6rkL9km5W+nSR5cm2k7C3pDUliWn8rXTLHcii60OMeaKR78Rc5f6gC
lm/zmdrFiO+gfKAfdXxJgMRovcZfgPI5TOMt3JNWcqYRPHJhaQMlnmlPKdjFa+Je
FdYqrop9TVcKgJ1rEd4JwNbaZ/j/REAdFbW+yIAk9sIbdS3/dIBchRONvpbpuoN9
Vo6C6xwuTA7nleBfGByr2lmFc+h3+0pQZ7vfrpn3xRLr7fN6vYG6criVIfmOCvIe
LVO0eaGMLBnrHESUDG3u8cCqcEBUaNZoiIec6+7A4+wQc/gcxKcQPrOAhg7IxcVT
ZV6zjjNGfQ/PAGsjn0/uyOvIYV0kwywoeH+Deaqbb/rr/ARZCC20v1l3uQvutvfo
fowT58w19CC/oKRDPqji5kKF1YhKO6BenkC6U6/MoIz13o9YwIn+0vuACuI3Q+yh
X7vqm1aTu5Llpg4P9uHWUAtkQXme3n2XJLaZIeoFo9tbsLLBAqKhdyBDrkzY1BgJ
vfrjs+ugxXqityiVxJ0YOy8UIL9P84qbSFfE2645/9FDBaUz64vy6/1xQsdRvFtT
X0CAhImkjX2AhKyPIDNvNtz5zT6ELfip0SEKbzOYQQsr9HxvYjPY3nHc9nhGWEgX
BppbsSfdoh8g3BrXodSB9SeitE/UroSN2jIK1RefQMgHHBjXC0Ze0bzGoulZb1bz
VogvBEoI/MUVgba2OMRUaXW9zYizCcm8Wy3CClDh5+omcSDNZV2L6g771/pbVMJh
1P+llSgGqnIMKl8v3w8zfaKMMS57RdbCAIiVQFIx9XdQHzW3dUe6K0l7C6QI9hYj
iPAHzKMC97Writ1CRWsnfTi6IUoo8I0hTeKZ+bjV7ijLZz0J764Q6OReiHbZa8ke
/vVnOpvJ5Tv7iy6xNwUNSHjvWrVTWx4mt93gn96Tj58lbZbXa2vXq4Oa0rbtVi4b
jOmjSAYIrU7alLoiZgLaUbwN/i+yJVsiSjULuNn78YGeIHdb/qN3AXezMFc8W0fF
YLpzkNyHi6dwqrjt9SjUZV7blyBUQGtuXnpKRurukRowQhdBqXrJ+9p6tGnUOz+f
dd1GOWPEqajHceA6oRZzwF+98FpUHtKrcDwb9D5V6lAlP3i/4kr8DeFDcyoPRYlp
cz3h/Oknp4IMSdeSij+vW8zunHmL4jJk34jM60CTWevlm26zUBYbOiQT+FB+tkUI
zhW+6S3PhR8uX89y/rLG7MZY1aHYI61Oei1YMiESgaJWQJrAOiMrOU/kP0L8JdYd
CSpajLws6A/r/EAeQ0JZ20kWSVqZqyHdQi+M9+yRKOT5fnBuKeGgfAx5dBC7/3xe
XYgHr/HMP5uxFec2Rkblef0Dwhy++F6/HHr30XQ2QZ9jQ8zMzQ3Fng7zAV9JtKiw
GB+nVXJja0E7jIkF8Jtnh2eVQyGQn4PIH+HmQ3/X2gC1GnElesyAVPkKTky13aBO
Dmej+V98Lr2AFTgZVPCmvBuaZo+vAciXnchPwkMRXlvwD3rSH1uQQC+yrmfYyRTU
OTV8m43dw2tBCabB6xPsFWt4zFX7yc3xlkKRHhJkMLWFuUdl7N9s1RbN2d7qjRd1
Gj0EhYwo7++SAX9K3icQTJs/kiwcIx5q6n06YDYI74XK9XhpVevTZrz5hzdmtOz2
RsrQc/eogj0BQ96WZPfX92XZOxsfA9jj+M2ZR4Xa0jnBNrAOy19tygM7KxXpCLuu
uZ3PwI0nykfFhEn2j3bzJQK7bJuUXJ3OA+IpkOQt64FPr3DWJExKfolZ2dkt4Xz9
m43FZSH2ewdF52+DFXWmZyHLgT6ReTYyjMOJpj6sYrTAdshLvs3bv/8SS2j/dzFX
eZ4stm7ctfWXRwVjE21iJYlt3OuaJ8bMkc9QAHojMaw7QOdOiuJRQo/MTbjVUdOZ
MlXTRTt+mv8s33Mq+ywQv0fLqyjn971nQ0tXzarxnAVvdFZsmo3vuQajT4swgkkP
ib4HLpPvC9QO5fzoJ8nk5Ue3UhaF4rRCrQWeNhquD/2SJPKaKH0PpP7i7dUEnjhq
b+32qB4GnEkp4ylRzUfcRdTQZ8nwJAxqDX6aI71vzyVLrNF0VDDXajzG0aVP/nwH
QmcqVLXu4O1H3SGrtT0TlAXLzLeSuPJ1BfqB7bU6dzojzaE8RKs4A8rmkAq3ihww
udSI4B+GFqbfmm+/VUHtAZpMCDbg6edq++DR5TIeqv+/QwR4ia9KK2rqljdlEj/S
ijFpE7UDHR4XblYsnpCpF210OJo5kjIpxP3LO6Jqy2fr+cqk75aEVW+Kqb3ocziJ
WrDo4+kLM4b9GIj88SmyasmpttAfZvmf+XVhi6wVOFaOfyLHB0FwUw25yNqwV+hs
ZsBFDalxiq+HLXHKI0G5ZMXMe47UeV0SOBvzTWLmmOT04CWlYnZgTef3EiBv7H1z
P5sVq9kBvViLHzUsfFp03o5s6y17QjPrhgrJ2HEz6K5HhdtkVvxS+QvQqOKgoOPN
y1/K6YtL9Nwq6wMjsEbcBCCkx0gd0AdbK2WyBQTEuOjp13aKSApSWMI1DuzB6AW2
zyoHxnsv+ifPMVnE0cj5rb/2tXQ0s9qTMHSoZN/WQiND9unGG3QjXK018kAGdqoG
Lll00NJ8Rbd/jaVuUVJWXdbyE5wDTk5/5MbwVDt3CbFUDLL+YAtm2izsET5QZn6w
xXgV3ir46Kh0tA/2XVneNAHWoh0jnfQsA86wIHITHa8horLEsORDKPfZikNgUwqs
2PbTkdmaJq617IeqI4+Ne6c9zmr//RNbOAhjuIXGZkb4uBcWogIagJL4a6upLHTj
y+X9OltvIafMaieuN717nsMAoLXT9JUxLqbmq3Vjb+ENROXG3hC/OkateEGr0V5M
50A9X3i96YIv5cfKCnHvEYE/Hu74Sf40UWwUP2rNeMT7qG5BUobm+pwAETMyllcz
8zEZppr0Wvcl3QyUdEgkC4QBQjvyEdnecv4nPn0OWfRphFAlcvL5lxhscDtgf/tH
QiSZ6E4bMgEBelwLfhIluRiJscdaVfAD8Kv7mMXHUcoaQuXMUgbVZwxVIuXryVfi
jxREmbpow1uz7t/qPczUQ/4qoH25VYowi2tV5dpe6m1M8PePNh45ThoDGYS1r7X7
s6AgD7D59LWISHCf3lASOkEEsyDt1REvfvfHO5v1guhtwTijFG9iCWvate9LGhoo
GiZSWoUyLeXq6KbOwqglNQZqGNOw7YIqmWa/zISyLOOfEJ9RGskDK7qd3QH/UTkG
ZhCYYUmjnIxuYZwEQOIz2Zq8mxlRcyAa+N9UVv5gXliWCfShBLrL6LjEDhiOV9kW
EXlaz5qUXbVFbChXnjIGhdHLPrT0atC8tiXg8xZgjzaPtxLtP/B43mYo4viAtxU7
rmkEq0tfR3Lrq1j3AAPEh6fVRDcwusDGbkA6NYfwWLvdSqXF04n/9EdyCTtoruX0
Pp3XnWhUbmnWOJreIxDKwi7NTxAqFi11wmThT4fPYYIkYn8UBHqEETuipexaTNj6
4hGIoczsrFtI9W5LA+TgNChRn/YkocmyhgMGTxR8QCjoMqYglGSY99j1JoBC/KYM
TKyfqM3qzCvABeMf9wMVwV/7/gi2Q3v+baybzgkx7io2vvcDQXEdZ5cW8L1vqnsb
9hwhhD5WcgFVF1zYoAOk+bAq38GjpxADJ/MWUEVu7qii7j5y3TFXNyjG5L7QhIPq
W8FJXPxqt3Vfq2tJLtAr/QNwf4JSwUGM+9cviHWQaxDI1sB4xJ/VBm6tVw7iwImQ
t95kk1IrcOgtEOiwkcycJpe1FrHyLkDu1PMfFIPYmTYT2HgXMDn4Xtbq2jbaYcJ/
8GUt58bbKkB4V+D4bokq+YmOnN/vPfGuYqE4k5cS99DZQRNlHeW9xcyERz3oCMPQ
dtYrkMDQqz2WEDCNEHsOfoxn1NaMBXrTOuzSYOYQ1/MIlpnlzGim9NRq1aySB6Vm
sO/xAoyQuvcgoIbw4DIRnhItHgBxtZIqz5qsWIGmCzlapEVSnW8HOUWFP3jkjweh
Zo+DsDpp99zNzVzdc1CKEvDZbSDokaoy7FX4zZmJcKA/r0R/j6lAUwzAys316BMM
Br+Wjt3GcSlgxIRfbZ7RyxQV2GPMcbPzM+b8sGhMTX/BF+uNtntuE2rT4jMt2lBZ
yBhOIyV0i5G1Ahv3nolZ5w778S7SRg6FdnBB+pHmJhDN7RBfZW1MLGp+DkXxYe7e
2iAPpvZbP/Yr+5/aXpij0Cavx21dSahkUV6Goz7sqKy8l3tbMtluYTxwwWX0PjbD
Am+LmlCeY97Bl91uoWJeKXB9TOTnVom9/vyttUIC+XFo648c+jkY/dr2dYT1wZ/D
XoN7I0peHHrgJ/21D7wtIyb0Ts7yJl6x/CxHEKpkvrcm4pGa0TXUYiS2u8qM7ZWF
0X3hcoV4kVAKWW9Hg1UhKtV9klHU3i5E7UjO27XjETWnGtwONP7UfhjMSCp9o0Fr
FYADX8KXPynfmPDEN6LSkaWZjcIexkAmyDZ7YHJgCQZROEHE+pnKYXG35YhfzmIY
lnYufV2sfKNBb2TePcKA911o1t0JuBvlbhHXC9duCallFq+WORJRtOkAVmPwb+tY
0AVe/vYbRsx45TZ7tM5ItaChfwGaNsknXffyJ8V/oMh19mhsL5J1VcnsQ4Xg1P/J
FBPj9g9z4gyf8J2LLUDHVEtpsitgO0oA7uXYdLG69XmJOaRJCF6WS6JrcEofyrhW
4MeVftGzpuPNlEMtk+jfeOu+klGIqwofLkLuno09mC1Id06IaCvbfXHwU8BbFOtL
KE2Bp6F5MWwt28X9V4oxvelXuT/3r5oz8Hdo43i1usMPstIOXqABPDVYkGC2Czk0
327KuliKmdQBBXlqLqoCcmnGHMT/Ee2anFp39FirhJm10K918hMMyShbJI0bHAHG
3mBHMNvBrMWEjPjroR0jnPG/lSF6SfjvTyONUatX4vDupvUjIdydWlAdI0ygkkJ9
nRyJm3Zvz3W0+UWwy1RpzauFhWI8azEHE83/AsujPhX/YKFLRatAPG0eW9c3M8Fi
dJtO26AvlDZH/5MBDdWyGZo/8R2XbtqQhgRtkQ9Ss8hvKQ3xlylxnHLMGwzn6iWu
Pdp89I1t2W50kLfu7RCYYcWr+sGKLcWETgStU5HqW8A3Nq3ZjIZYZmPivW8foZsk
tIOJLfFZeq1OkkT6QpWxKyPdAQoel05pEpJseRRrRfPq52PUpQC1Bhhv5WUqEZOj
v3zyMI8mWsgMqQ9Mq3YonfTry9TZpCmvFCGcFSiMTeKxCK8PpJ/fCNARwljl06HS
b6lGyD9hK8CqP6rUh1INvyuE2m0bDO2/+IX+MJWv/huOfBeq3Dk5xLrTYJ7RCDYi
yeTjlfUCWqd8bLdmATu+vjJlLA5Hd/qj67deRi4Vbho=
`pragma protect end_protected

// Copyright (C) 2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std
// ALTERA_TIMESTAMP:Thu Sep 13 06:32:41 PDT 2018
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
DED5BbxcLCrzgr2tytGZTX8Rkov9BImleRk4E0h7G60qQ+NTDEYQaNi/Ogua937I
bzZSDr+rXASKQ2nDQqQI5hFUSiNzD4ryuIrDwHf8Q9rBrmR2Q8V2QR0BuheQntVn
6EtE929Q8sA+hixGpumJb9n35JMsPui9+6GSG3KTN7I=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 18352)
SnwvsLDAi0/ILVuNCyjilHVNA0uMp5U3APymBVrwfhMipOVOUBaiz92EXGx8UZDI
IWnwVWomfVhxS1rcuMOBFATMgVszfPyLKueqQ3AMsFq57Clp4GezYDa1qgwvo1/p
5Ou8BzcBroD+fmicocdvQWgjCA5HH35XLsavJpm6Br/wXmuJRygD12oHXXuU8bnK
KCwIXZUMowCAkk3hepyZYul/+lvAfmJfdDN3/5WFpywBtnbs1CI8VWqOoql1jGPx
W7VkS7yQ/Zz0yItDptI7ErV0or4A3rPRQreDqnVtgmA3Xo4214kOiFTt/oNqkWP0
RWIlzfeQJ9twRvufuYtTLZbGRyzWBOLupKeZBqWDjsJ3wA6lkanmhANy2ihzziZs
ObM90VZOMwl5LLbzvj3HAwq5SmwR6EwdSwgcbLH0FBZNsJ2lUX6w28yr9xl2DImR
fHMS1neYhD2MzBKKTMclbHxyKrNuiJ4uP4oj9GmraDtJfmRATnQ1IVS2WLZGJoIY
CTVujU8He+cLDGL0Zd8eSTg+q5ab3Ft9072cehXEL1IHMJFhfA5BQDEi8ovOhv+9
f2sGJa5PwC2T4WJ+No07KbSpoUVxoGNpRfOZGWJ2D7hpG1udV4RwVG26YGQWr/Wh
pGSLHLpBmEv6f9If7QpZ+DtPt+nSYhwmdPNEVwd+NrJV1JkjZDBRJ3Bg3jgPMSpt
l0DzJHJA//188SygLMbAfSeoMIh/JKkMM0NaEj/lF9WJ25Xts0flx8x2Vv8d/S7+
SjH+tm2iPyOIIJYAoB+8jWDt9l6vDK9TQoiO3QQDojfu1zNFkqYcU1P8xQGbTuVC
2JzYWt43V4WVDm14UXJZzEwBDKNlPaUbV8R3C0evqFO+Z0A9aO9gvzG9Wcc/470L
PHnCLv2IU/45etgHz04ZbgRIQ1KViGKMIYN/GV1TAVZ48H1X/ICEVImXDJyKrkiw
j8mBy7qZ6bDxPqBw0cCnLJ8XtCeifSsa1Xv01gNbyOC/J9R4Jidr2WQnyxx3CbKc
A6Pd/Hdjc8AN1U1DWAJvll/kRFHgHiCaJg/SEJCRa9z6E/SlOdLdaowMzGdAmwBb
qgbHNuG+HWeleTWvKUANI6UCv556m7kBXXjs1pPM6ojxmGcUDviFjAKPLWoWaTyd
WzYN9QRg3qtWUmDYc/Rr8LdrLAkZIChmBtCH75WDTlDiotrxyFhGLHiiPpidxFqr
Lx8g5VJVLs3vCrAlqkOJvVDVUGnJe983HtjkinmLIqryiZAis+EyByGSgzcHmBip
+FXizAmx+y5Zbw7HNZFCvrwHP+dVDsNTjVEHbaYIRYnPGRcKFgAe4NLFrcU8oCN2
sa6TzROMVMC3MNbgkXFiIqwRyHiNR1eV7LVsiV0S/8EG3ROQpkmgTch8MJreMWha
6ySEKSB7WwK92eTCsvGT41ullhfnvsE6bFZhezy4sxtsiYv89hPFaq7QJK5OGtbQ
3ywy2fzKUWf7YJsbbgRDxPIyqpw6FE3ABTFu6pxUar8Mr5JWGlEb783KMvzFrTcU
fL+pkNqsdZZrvx4HUH2xkOgCyIe6xit7yfwvryPZNym3SEMkoSjDEER2mv7KxQmY
+C7aEvVEfJrD94njyyoadQA9X0Nk+lBPUkldDcFL3rdvQ3L972fHJXf09NE4kRPz
7MgwxUH4JuFwBg7yimrqyyY+YqUuWntKSBAX5Qjx0xLawPYUpw5gs7fz4jHsF2TX
QWxEQUgrGIkJksmUzzu7nBf2rS/3ZUPCB04dLS70y/wlDsLrps9ttiADmZ8fu9k7
i9y2aesGKp5L2ENJxsQ8EuM/l82m0h908Vgoh8BRh8pGLZGFkYo+N3hndIb4NaYU
BAPk6gRToAwmB1mRLtOQ8sI1BcQAaCELfZuPwi3esMFlLolVocZ5udiVSS//w8x4
tM9HSZMYAIDLfJGBwf4URnDQ18mikQd6JNTIRA92w4JlL7gKzW5o0bdycWEgek5N
gMZYlOv115gdKDmwnCZKXuISCWSXLgHRjPnHpghXTh+5pruglHamXCVVXTmsW4+e
QZmRE7zYBZaepmN9Xv11EoRgkgtkIr56zYko754IljGUpAzWa4+h9kEIZOk+78Tl
yzsKbqxw6Ymv7/9wt5JVHTMxDAL2HJganeZ5ch9r8lVWdymMZQgja5QkHz8Nsw/h
6Ybvlz4Gk1fd+vlffjlKZMm5KVO9yG+pDzFiMkmyQx8YelWGgn4Xs9V9GqaueQwS
+vKmZJ8PoAlDDX0g/aTklFP+uLSfADJraxhKZi/qIfa3U5qHRZLoHd+Pctzm8YTQ
EL1soJ77IODIb7qXG6Ubs0aX7UmkW+mYDuwnbLURfLGzVRSnnPjdAPdLl3gbyhKa
z2PIWRww+uR4yMAnxMZO2xVc3unLDvV7L2h48Wh1ScbX/g4lC3a7Y50BmIlX9J8h
McKvVFGvKp2UKf62f83AtlnizsAAt839iZR+0kIcSu916ueiUei3+Zh6/JPO6pJG
rL0Y4JvSI+eQ7SkBvrCHjerB89j0tgTZ2F8ZyDHlVqMp2j2gkXOI/ZxHMB13X/Jv
2kkTyHkaHFoXUTxKYah1ZEOiLlN3pBstzWLufnjLclcSv3KzU9RHPC1jwvSkqhM4
i4HKeWHkFfV4J4SN+fJrCwJPzcFqh1klGdvyTDXQCpab65Q8OQ0REcdqP25U9ZJ7
lhSOklgMQ6mGgFYaquyW152MJOrdcGJKmxO16d7/E2L/OgGEmwyudYvTMxq0EHTY
kPe97rnEmtKbvjP2T0TForwlHmMvgkp1Q6planG1115VmgCnF1+oEk35wBwXVK7o
NyApFVY1pCUzsZfzei8wcY5WARGGNALAOS8rnmdcH6lOKkBy3S2Ni7RhKFdnQ+zd
f8ON6UW+4JFHA9b4GXeWMqDCHhp8mzaB2yfIZrc5/hPvdHcc+SBOU8wQmiodT8zK
45eRw//8GYw50HB/mQTOqMZFmAahjK+8AAvrQ+EfdnXRGLtNF1qKe7auP0CX4V+a
RvWAv3wqAps60F4FkglLAFLozfk2+m11zMJ/k7h7c5ut+fsgd5AYuBbJ8UQmoreU
8GgJ/BHc/ZSoHkIWnXXvtGyBdUbhxOfvar6mMJMMN4L/FmabLGpUJCyBOq5lqqKt
uX1cbBDZ1UwCxwjeandteU4DJ7j9CpKHRneX6yBtXkDnfawAsLLZg8WRtSGhrNcS
Yf6uuTc7fEjvas84XMfZJH9QUWqaQeoHNDLb4GBEIguQNcdZGHknebz3QsjSb5Ls
SzWGVSnPZipcAbVlzhilCDDMB8h4MEzUMlLOYSvQeCLz6q3h0AFz7nVVW+wULBxk
J898W9vAY+kO7uYEHaLkDKkZpYd+hpMc7IMqwesef6Jyuer2X2Ge84F6288R9VTn
Bs6RCm86kcZ49j5gK2c5T4AQ4fs4Q9uhffD/ObGQT2ulIoOhqSmU8rHZ5TQapGR9
c7JkB0oPuPt0KEEVPctFKBwdvgDC/peUDVcf9CeazwQ4NbjSeVZVy+OHlCjJBC26
V3DqoztR8gIY8Q0a4S8hIVKMcDT3U+SzWa2ER67xK6+ykSJqYVheKFUhXFHNsskf
KvYOeej3o8/du848osMbnVfA3qnfqDRW7j5IHZ4/++5sZQePMwysQz1Hj2ikejHc
WVh40wWrVaaExRPs5srzOH3hkl8jVV2FKYmKlBvBQkE7os01ygOAegtmi1SZHgDv
5IDxrnLWU0UUHDgwBX7A+JspE0lh/C3AOcDC5+lXdBqwr6PUdNQtW1fB33jNHt1R
MFw8SVMexbUiBaeSCh/3geAK4uFRb213d0HkqZ2Fdjolj2gEQOYn5moJqhMikftm
FIc6NiGKl/jYZ3q4C/d7+An216TC5eeN0QtYt8UyxlHabeFqbaapINbmP336cNTx
U9Mr8yP20flqWO1SWBHsjSoGmNgzDR2XsnO7C+c2dTUIrv5OcQdODDqwcBaWyUOQ
7E/JUl5979LPKg6ZXIU+Y6CvQ3sqmswUlL8mXM+aA5AxdHiaDpqB9cJ5UL4D8xCE
meWikEaFIDh5+7JPiKlbiFNnTYedJIks2oabJjCriB1OsbASRYGGVUM9gWYfZd9k
fkYVFCYOVd+HiUUxVE5bgVgvzL225fdlzRDLzZ8F+nLJix2k8DKpKG1KzVdb89jJ
IJbU4yuPMo9oK91mXCfaaUS/THgiMluDzjw1+j7K3B8j58xFvSHPpZKoB8ok30eS
KAas7vZQNCeEWY/YR5lFkJIhZbtTiwECmeX5svccKkCnIm90yZB1KEkxrIotnET/
K1fDaKtF4Gn9T94eoo5URgAZfaQyZf7zBMxL8BVP1exhpT3nts5Mqh/8bjJzi0ZJ
uHKcvMd7PK+UWdhJwPHIab6Kc7eys+4FjNHKJsXqznyzd1UKSj8E/jlAUK5fubXj
cuelgl6fnUyN4hwCRFPfXxG38bxr0ZAWIrPvJ+tixa+yHxIi7AAj6dmIVUcWAXTO
JcaNMYTPM2eWEAyfqJpeaZ1u9p793yTr1ABL+HUmIL12FJJ9Jn7F97t1Nz5BnSSz
PIVWmQlqmpRt+E8zsfAwy/LNvF2DW0y5F/EGAR4MqceqScsZg/3N4Cm/ZHYz9HL3
XC+u677F2MWR9lIviHaA8iDNRo1MbXwST7rxNSeoZ6YO001DnnYRUAzMhsGFcmOw
8aCml+9lXC2FyQhvO1GIlrWUPN0kgxn8jeZ8kFl+CfVAekJDmK1KNUa7UHlH/Vr1
yNXKQWuKyZN2nrP3L4wGpD+Dm6NJOLo3vgQgsFRVEA5X07RirSau61fFy17XknE0
zMElyKEMrmrTl+Z0BTgr07gAgXcOjPXzF0Rycg0Oo/BpMoSCtiKX/vGxO4XSG3Ud
8sziy0C3ZABNcjC4BhmGlXMKbiiBPoWglcrtRQ6pGJBgSK8VdUTj8MvZpcwakMrl
zyExIypEnxD+6sp/CHg522kCc+iew+HydYUTm1wa0antpGu18NCf9qgvwlfrgm8K
XRZaB3j5KOZAIS3QVT5j9QaLgvQBtPFkxVUwkB+rTGcukJadkyWh9aItb6zyegN0
HPAn9p1w2LS/dPDtCYth5JxsjjLlZ3fwSRcXoxCjE3RjynFeTWj33do/FKW8PLZ/
kzPH75xy/hTs7veHvAkaxO+Qm4zLx3y9ndJG/QYjyzxJeEraSbFHudTjeW50g7Aq
o3b0mNRwOxZAvjnHJDrdwH/xNr+qA1WVBsXjNAGsblhKXmKWVZhmY4Fe6YSEjVLc
ysGJQXdf+5a6gxkqoObrIzA6H+DRgmvrCWi7ql7CRsbBjLevxCpA2F1RrVXnRUqb
aWVfn3a/WkKB1BDGgt1z7z7UrjFHAUrZSi18+lMuqNG6zlDLxZD0uEaYh14xqbcv
NIv++ONbHVKQ/AWgkfyIlBSkJH48KlrKXjCgqogUX3NcIkDB3zzxSsIZnIsJou3D
R4bqj/PauFG+BVq25dVLeNkZSIMr8C7wTl5sQEcg/LVyTPtMvjREnmS5KN+5yq2Y
2tF46nApazIoV22sF0xjYCU8FXUgrzu2vx4JhqGh3dKl7mmYitK/3bRx8c7Momj/
wlQp6UI0J2iekkFbS4YStbSJnDR/R1Rlc6GRTnRHTEg2N49Py8AYPVBPT19Ug+Eu
JK5uVBJk61szuP/eThw5bLHgDBjn5rjxiauykiimRX5LutC4Eeapq27XL0o4Vwt2
SUBIwMRSJB61m+hSm6VZAx971ZCx+n79IZw29tN+/0bLn3iTJ4SnmAxXuwPSYVHH
U9usEst5XvUZZyxU+kkhlLF2F/sjwxvW0mVTeHljqq6WNA/3eZc3+lyxkhvINhd3
5AaKUMT2DadWhq0i3ainBSgbTNIm6E9HPk/PCY5sSRlpQT54cnX2i6/PTpN8TfI+
VVzerELBs0PA2t9oxBeGAc/+YlGRCsidFeRdlSGWxTOJ2JyYuec760SJDNN+tbLn
uW7Iq2O6zw9G46TZvGvBhSIngdLd0dkfGo6c7JL2+dv4XecBbqplsFa0D+8BQ5It
uWuDZMuPByNf6LYHPza+XbseGz4KRl3nSyc3zSK5l3RD/H77KQALI86mH1flMGIA
PLsi+iaajuUf/AQWrnB1Zb8GdtybW8bQbb9NZcJUYEsjBAFbPO1CpTOgG//4ZXMJ
Den/k9VMnGeK8QvKuUClpvV39WamEkJVJSrYkOl8Fbqzll/k3zea0caYM61WEw+V
SYEQJzfAMmcELTiSibtK0diX1foOMcSy4S4dpgrbT6nuQr4uq8/lS+DqTlmHcaa7
HX1iq63yxNjmANpQrZXh01FqsRDSo7auHyPqHBLvRcy2k8Ks+F/zYvalyPZKv6Be
7KxUkCoyzy7veqL2DJfr9TWPD8NDr26HwfLnegfR+db+ml6/ojOl1jfDgfJ51m7j
Pb9PUBiE20vepfq8E/KK/dh/O5QC1m/NKSTq8bX7Wd1pBDRtGpVFMujiJ4pLki0r
4BE9pR8o7DDXXAhQi4YC3sLS8uRhUxZubuxwz2pOa/tVj7RyEVy0ZigPMoEjA286
6UUiwdmHn1OBSmTzzj4v7CQquvkMgXtM33rBCTatMC0Hr6B4DYS2SBPFhyAIQz3M
i5MAt3iACJodKPlVKYCtD3J+H+O/4Q44QpCIn9eEjqyS7x6lHvtOGibv8NmME6RZ
lMSv7NwFXn5dHipEdHzYvuZVrczNq1ANZdODPhs8cmL0X+aR4FzRQ8GiacrvVFIR
b1y9ekNummf8/6eCCdT3ZmTCSTh+RXnee2/gmEDfCllPXzmkvGGLptPXfWUFkxps
MwsOX90qCieg9exIpLR/Zn0mwzEjcRB0xIgToF7inoLFhiCszKD3QiL/OSfuPqZ4
iZMBXaD4laecYkOhq8oGXXg+hVFS/DQykzKLvze7Zj7q/i+6k7n5Enn2p0I4hA6k
cmZ9aVh0mpvyzwMPCUtSIKiLkJyaiB+zSD9kZPcL9V8MHGw+3kErb1+bwSr7whe6
blphGp3le1l6Xblm/JkrnEamr0jrkGrjm9YjI9QQJ68JyL4QF4xzPhtGoXFnnlNZ
kcN2V6uaYbHsiGV758q47LJhatMZ6XohWhxRoXXCA2MZeDtqYFld6Rbe1325hLrs
WtHdGRKh19+8CqyUwLT44oDXVj/u+A1W4V3XDZuhyBWX3WikcaTNuv6qpLvZuxHC
2trr4A1vE0mvqGLsgkjEUpGsuhgcqD+m2ntzg0MJPHcJ3RXdKO6Kugfy65n+zvm0
GlwM/Aib4PxkRFUG7mFMovnMAh7iiIRXQvwflMgf29rbSaDYSyF2wgqFshSREVde
tBMD+aBfXeIyM8o1ezGsURIlcWdsF/YdRnWwkdhH0opV26xPK78Laet6gc1SufsV
LtEul0hzJ86ITV2uPtos9EYgExT54WN5X+/+r3fMMHQw7kpN8qFN3FBD9xyeYPuh
HMVkzRxSEDT4S8QJKAHTgySJ6UWdXPjDuQ9PJeWKCgMJIcgKx94qfsj7Or0AU7w1
B5H9oL2swF3qKZjZ7J427nwb0CquIOMxx3N9/23uoE4RZ3ZRdKAG+Bl6RcXDRqeB
RSfCogjzPKNseh8bSvtiauxjcnv0mROxXXAO6Mmq6kf8XBkTnZAPFZiTXzOtjKtV
zdUMxHIF71aENtghSxbqOh/1+4FIm2N5h13nqsAhbr3VUQmSHuNByDwqxD8HOON1
zAMif7aLqjSeFfTo3ihVCUH/F+8UABbGJ55NVwTXBblxbALQEUxkdXpn5Bs255wJ
yIRBP6szx/5EVP+IN92NT4OdRm43QPHOvNvsHIv2mrIU75P1GT0sr4gk4ae58dzQ
/SKDGNKsGP9QDfQ83SnZm7AjG4PCb/Ycp3nn4pZLQmUsWAZjz29t/bj76X4nxviv
Z/W4X06/pOcO2RJ+wZAWgfkfXr7eUoNlZMXZCHHPiGSU8P1bFRXc+U0zNGF9dIvb
pPjlVMqugnAcvDApyXCVME5/sAOUntR3T6/bQX5+WJLJH2cWna8NBV5iJnCYHVLP
K/IYQbhgEN/i6KB/fc+F/DkxJKRBOK8PRAN+EaRTb0OuMRRT/96tdvhh9n6MRgq2
d209wXP/OXzovGFCLhhH4ZZdcPpOsnl6eUyXBo2zmIdKXewCVaz8ibTMZ+g95fgm
d47JjvIFu3Bn4I9Z/mLr2a8JXE6E4jvrXolt8fYAHYRyIjikSjFLbwii0mm0H/bV
uOHqGknOtSEu8R7jaPHYFUfQgKJ2of2NfykSmnO0cHhAtmAE0GCa5UsDyWlXmh8M
D0M9R9FyAoTyJswm7MWj0DZh7cc8kYZA2CFNE/i8ffPlMguuq22goy/wWs8Zzhql
zGWQLNaiksvp7pygiKHshFUXJzdJjoNZXCDVd2ULdsEww5OejHN4hzyRaOzBcJxZ
cx/ulpCdiHzCoE+2LxZT8C2Gd+mTvNZIpEqW1HAWVECCyO6E7BqtPaoWbDnuUi32
0gLjyx18C5ubUuDNK9+HBAx4VluD0sl1/zZ9zjx7Qmjemv89/hoJEHthmxZ5wqUE
4GXjkHR4jp4wfWB6jNrYvOMQte6cVyI27sEOun6oXCB8YRjvCe3CI/q52gEJS1OI
+hjjqGj8neVowhNnPXcu/UuWTifHxx2/njB7LUBmifzxkh0fq9nnBMkThvl+J+vy
lGKJSNTHs2QdCef7JayTTZ4BKkt2RzLS/0TJfQavSjOLvnPnQjqGEVHretIcXgw4
1QGjXfMZNkpgzz21vTVrcG2ef8GjsOk/8rjn5hkZsX6j9zAHkbr20zxpsJA390ba
bEdGzL5nkODdwclUWvazeI3RJlH/T2aiWJJUi/0+OIlolaDNnxtP3H9BnBgxlxLM
0TDGFHw8l3ifj5OqhZRr+FYRo4AadGjxhPqb/J3CCwWc8ktToJC3faxZHeimxUT2
LsY59JihUUBz8NIyYm4WKpThmRm61Fpo02/GEqsNhdEUi4Myz28O3fakI5T9/8fW
xpVA7N6fiE+Fh6fpoPgNYEbbgdwRlEY83jhjTVjmvSl5SkFJtsZXB09agXQFitY6
ZiwN4Ji0e+VEZ3Oxj+VVPN2ymp5wX01YUGb5xEDHPEvgbmzXH0L1A16YW+ddTd/y
JkFWQw7Ep9DHa6b2v3Anwo6C6dPegCZrF/+L9MOBLldqxO2d5HwkFNuQXliHFYPh
UsGMHqecixp7fyrRkhFVK8EMdHE24oi2wAlZNjj6xyvmtMh0JQTrsT/rtOLH966v
5gi/L/R5i3WEhLL/sNFjI7WzCQb40IxDMB9I1YXxYIJWaLxQIbEiExrmGsDdq9F7
+5wGPzwhrbpbXXE9boazqGQDs5NBBs1LinyPJFc83ATKRbznrOqEKaesEu4IGEIC
DoSKfO5cfXQEjugQsgJEjUUK2OgC6O2fIgB+DKaa8HUcMz6XWxJMK+L73E/dfMxh
Hs3+uxuXmybXxzu8WuSBTjS7y8ED0Kw9f1f6qT5vyxhKW1KILc6TBTuycrBGVE7c
3BwBWimFGgpKKMjU0WsBSEm6KIMZKE8pWpuwSu3S4sdey+cC61StsDu1JhLP5xKb
LYf1jpxwaSBTnZ2Iq0NcjDogizHg3eHisyYLC/LiTu8SJn9K0JKqq+aNsVyWu7H4
Hy2qXOJU8hflQIzVFH9MJEYjyKX6gbKKIaTlZtVRdJ+hOvjEOb66IYWuvB6bpfEm
pI3jgZ9LQHRgyFEwupMP5BTGdCV97PklUkk6hCgxpSP9vTUDon7/CZUF1Ike4aDm
hCQab2VNZqZtplkA6rL76BHxpWM7eHNzwoLHjWq6yDTx95H/XfGG4ppJDM9lkm43
JyrUHEujq66IGzVElA4YHze4dVyEU2mFc+W4Hl6g4YeioqtplGTJpA1ZXOHaQ3Es
O4L86Vz5nKZCdxq0Kjf1JlEJjg8Vj0aGGTdPm4R6z5r5KanCyYgYyF5+Nr2KQ4N7
Yc6YKxy3h2F7NAKXGEztx4txBMckAQtSlNiiAgjA/OD6WVjkMFmv+dAeMfXjUo+s
4a6GZZNV4WzVxGZhEL0oXxeXg4fAVvbDdd27qs2FZCGuGlYDQbg67f7/TfETOhGS
mXddJ0xt6Aj8xl4rs+pIFFIjacfNHmmus/mcbxeD+NF6QeiZ8EKYiDJRbJMQmeYx
rPyQLpJLNCLMrKDDYYVDINjYU+3wCC3+gU3L21VcoxMHjf0TTZ5X9a1mLxwzzU62
O5beJzbHbvRZkcF3Whj374PAtt+L1fIng7AWWLxk0B68mUjiwUBSI+APnDBSeDnp
zQ3JK527CZvJC2qYuxLxfJes2ouOmyHs38yiQYLLHLHuV3coSXf5Ew7OFgefqW7P
xhXhH7ffVz+Y6P+Yz13D2Xrd1ZQDcyUr6kLCAKoF+Icqw8gKnRW5w+BELdgxZ8xy
LJ19zQL7nMUooRw08rLMGnk1vM6gx5UnPi3XkbcUVsDubWMEqGJa5Ka9ayh7vSDR
w1YS5SAdrl8KzC1mynirNFYgvjA3qQ+6UEpvrWpXRCr/APWhLKKo971mRUWrq8MU
CSSVt+30GC27JuTIkDcQ3RLuX8MSSFT8c9odN8BzzBjDOMvF7aGL1jmfslOM9BqC
WlGPt0wbiIQ90Q3Lpp0cYI1vB+vJ9NrF5gTqzqF3rITbvtmmeR3ROZbqK0HGSx2h
FLqztSvwx1al0+2f9nCuxhtGMjwtpgH5BA1KdRgtpcyWDMGW/Q3m0FL9JCbcIqFq
VWiZrAqE4BDLW3JIczjbR3VacWOCzArigT4CkGetenGKi9LLeyVKohodiMZ3nnM0
v6wks5T+/a5X9GdOhU4Xs2KZXs3RpmD9RCsvMqy8Xqjrn3QUDBWXz5jQsiSjbUWC
tu1MiRx2ss9x2FpRSumZJxgJp0Y2Sn8h3MCZVjPMdATQ0rLmTTofl8iPK7BygIoL
Ba/yBw9TqEfZtALgL+h3OezGF2Z+NXVEmDgSOQwFSfwpzrdO9ZDrcPuVzOuLulML
O7gg2X/kzRCJ3dPPu4PdmDnmkJnl/SIZv2dwWU0jD6Gk/+tqOgNoVKjRWBwFfbC9
ElAtWSfL9+RiOjTlVBbq0066S1mh3TSE+Qnr1zD/S8iJcL6j5+cV9Hqx7AOPc05h
ZcbpQHgXUZjspHmE/IcsPRSJrUol05AQCfm9B5vkdM7FAk3T2LRdf38r6izA5hfp
dR90LFQzeV5slmE1EjLSjNB1BQ7rPvaCl16UQ9mBSrrMS3OZXqPcwiLlK3ViUgXb
6meO7OJBbHAxryT0zDCApFhkFLXbtzai4rmB4d2OmcmK9LrZXIsob2OZZ9Hxuq2j
aFHhq0K/hDxfUl/mBNwzm9hDl1H/hYh8DE6TCwb2elUWAZMZk1XCvgF36Vcwkh7J
L5UIDT5sxrKcov8Kj7HgoaF5QtDCi4lqTqsnytijg906qGSqb+rrMbxmIoaYGws3
smSLd9QoxWvYk8Q3j8dhkXLjwvXkxKt6aCgEOr/uX7pcwXbdtQPhMg3JfdBg/Vhn
P6IEi2EOxnWg9cCVMdtNA2BOuPC+Nqup4bEKqsVFcWEGm5BVvtF/InwtqAERYqeB
l5VXLNmHZj4I7XrOh1s98r6zpzJQ3iVav9agiu7YahKPkaS/CCCgeSEbM6a516iS
1Fv4sjGVD+JUz5jBTI9mjytDdQK57d2zvmXKfahxUUe6OQaAgryYvLzHLDCWYzoA
nkVOaFwWM2brLiaP9Q+cd8BUEG8LPetiuGjPiVjVJqSOulpcKxsAmLLJR5nQV9+q
fGyoCwGpnPjGXQuL9iYA7IK3M7UCQqw7/B6F1IGcRty+CweKuz9RIjwDKmdUiW1K
mSps8xjrP6aycCmUV+g8cbpabufeqD8LX7LKMkc8ZrlJU8U5qMG5qBlZZfXEPQP/
NJJsXxWKXxSguUlelOG/9z5+k7r42oyEUt9hHm7OYyg6AyslDbEP0qFh+oIKwE49
VAFLXgAAkvCACIOmUZqbm+m4mWkFEvlmZH2L49U1KvtF62IXGEzpTbmkCz+sR9Le
xm5amvnMjStXuVlCndHkXmOnnt3VRxPB8x8KO7W+da+YvhT1RSCXrn6R/hl+k5Ss
TQv3C+KVcS9zWSvR2Eb1cyiZRGyIpLsCUQSzxTCylDuOcHQPlapnX4MrBPCkF3q/
d/EwgZlneynKlRNtc4r0kyAj2vRfz0L475N/JQnB8ruhpnTOjdd3nmoEtfEitZGi
ls1PpA0g7hsD8cNJlvJclUQVeNvtWQKJB69D9nHyjq6zGoPik++EWsCFRAcXtTbG
4N+2PHiXroBXv7LHg1PebPY2YVXy0ZL6NA8A3QMruA9YYn56P9sZWY7V5GFJUFB1
ClogwyuI1Ug7d03BiRXlAyz8Yxumljdf5x5MrHrY4dpF35+j3O6NCOTr2w4DAbUk
Ohu4tuRj9yFnErAVKPDmaQcKR1aNXdXMkkRbHT7wLZ7nPvnbQlpVm4ABOWxniTGN
YaFE+ZZzk81yNlHQt3m+UCFTWHSghPiE4EwqqQKx+t1w3QYjDIfcHwWqLHab4XCt
xDxS1ZhOkZ3u5za905ahRzBCuZP0ppt2olFwxzp4mDjnKDpZRkqvZ9kFmvLy33h9
s/HCG+FJwDW1mw6qgfLSUgz7DWqg+hu391/xJAX+3uiEksKh+UvQFUX+5sd6FAf5
/9uWfhOzsWQmLusTSDIeoIVPfMaUgbfSANwKrmgfzP7Jvdm/KTcdojVoK3YBxNbj
d3tkP26asfovtlUZmgRij7cJkuBAL6YEAfe0H1oUua6qmMUPj1sBNDzKjSXIZEJn
tukFtZIH1oeY7hhPWG/b+QoaZg5+Fs/DyTlFLNl6tsxf3c1JXAhfSkrcu9Nv7tWJ
TzuRNp0Oy1iXD0n5Vm30ZUSogdmzeClKfjoduR8gT52UcmDDNW8nOCy83HMSgkcT
+RZ9sZ1dFltyCR9yV1wRaAQMJGS1w4HJ5XtwHAQtzfpxqJxCdOFFLZGHIqjDrcws
T0tTrXL5r0VbBrgUzBhVR5+pnWQa4ieiJjlX1y0JVybtEYD25jiJDV3/K+7oTPxn
gL33TUFpB2ZJBPPkRwAfFO8eaf48/t3giDEedMSPxR8K5PFSJRTaIjkehvSW2AIs
5WACnXIHGqMe4fpKoWE/cYeMzi0fpu1zOrmyI+twiC6bsp0At5vb67hIb7xBMsgb
kOLUwvmI+xlyOwPY7bPgh5Mku8Z+cHChkpZkMGoDXf1yiVqtbnVDXk4eSJ1ZDLZX
9mECTvbU8q6RbzhYiNJXwYXBNN1CSwrZWDAGI3frE6aq/zTRbvRRlEFfsZ8jsXi5
6mSGB5Nm8MitgXMEzV1ynxP6pgyRxe8lrhSvZdmEk2fb00q480Ic/DeLt4j98oHQ
9VuTKmGp96gfZzwM2V+L5LcPOSsN6XzVwh+XqYYOteefbfi77CxNRBJdSHcPmEXK
/hkLKpkWTYZmH+nW+nJxNyIoOYerqbwBPkf9Ov7a1ZekDk9A+g5nuVDwQ1Tte5Ih
+1bPsuIczGtgmb8JmBTlTdIoB0ckVX/EVuDtjBEhl4xIgn7y3HaNbq4VJbGju+cz
xgeC7ASiSYq6ie8YLIqaVlKunsq1+Wz3Ffk0MnKQNGpz4gffCyEJagjV9GaFFVQW
fIbvjN6TNKS5oTK66AoPQ6xn4lt5b5eb8/OGY3pG4agC1C5a4N3SYt4ZtmJC1hus
iz9lMwdqg1GOv5F8uDpYCKc9MG56CwSVCRx+g2FcrvlqlUjEKUee3oeTlaCgBHi5
QwhCrw+0r3yOJAikxEtAx4PCicinvDgpjedr/USZunTDr91IGanQBBr6Ztf8OLCR
nZKKSWW7CfP1uFG+Z6Zznytvco8G7SExMyf0AGBdAFuqXbFqoJ/mC2paKQebMvr8
BG+uA1GD0iE71VThNfugAeWIFFA87UhQWDEFzeo46Mkj7J/GM3XQUja2Ru2fqaHq
dzhosDIbVHDab3WG1/Gl90ELueNaoNZT/cwbqSVQ1aN/DwTtcSb0gpVZgk4zO0qR
e+T09MdbKKi3eZiVmlzmdvom3bA14dLBGQAabpk2iZ5gZp1Dq8VZ2v9jIC6j3szu
xU2J2VG/1+WoygR/FffuFb/DfP4ED+gN1Ypw64VU1u1BFgW8AX4CnXxH4xwzvvgz
FwalkwKM8Cw8sJDmz2j2P+RLCjpXaRPoBVpNGpJT2HSdP+WG8g/6APRsUVDU8C0I
BaE/bykmiePzKPPPDecXnI+2MyXOMvlwWaXQjCqRU4+WltJhdpiibA9RqKjXcxKS
zduBp5mHwQ2TpVKBYr0s3NGu+wCqBxR0kMFj0QELYz8CPsYT++VUMRgcAqpYWXxc
8w2Oj5EWYtne1oglCM8kl+UewaNSz3ZWd1MaXWj+rwouC8/ThxFVJkjrzGe/x0kU
A1YU4ZfXHJtG3EUWAEoHtHa0EndBItoXK45V451ghrIeLbBsAD6NERW3EO1Yh0If
etpG+fNyrr+dGCHzlbsgpik3AKmsZyoaSgplrNO6NBL03g2rKHyfmjfSJoTSSEZ7
7Ww+tqRPA3dc0w58/dTnWeSrRkivaqSEjMmApnyrgkTYqS/p1cckFQfA1l72Re6h
fkPG/Y1A+hyNH1jrTH2i2D1SSt/HHm/7veUg8tvr/eJ4tCV/5XxwLVY7Jeu0jhTX
iv6xnIVvXXLpKCLwgYOslLXfzsEx1AjoxPyvFBtahr68k/pdkj1HUSntIOts4q7l
oc2m9e7m1y4qdv89OuPMl12yHG63kiW2Dnp6nOPjYNwRDgQQVwKKY+sZGIOK9r97
IB/m3uIgi5m8n3SMqdPhqtRQ/gErlRn/feARKipFSWQHHrV61V9H5up8Jd93P82u
g2SlGiwFmmffR9dVRfb3tzR3GKrXZQIIc4VpTxzFok9z1giZ9n9ZNMpglgakkHG5
9BMLvEXApf7DG9iVoP9i5DhYKFu5VMmYge821iFa3LcP8MWPZRFDll9fsL67CVV6
XP0JtEjhQhCvDmcY3KJS/aBJlJaCL2F5Np9cM4kH7V+hLlKj7LlZkpByIBEw0HRT
qZ83lswgMdU5qGVOZeasKBtALTL8n9oMbc+jaQrBv8WQH+lkNvt0RqqxbqmLXVO4
Y9ex+4cEFdv4jnGU3ljXYWo2v/HPjy+6y2bE0658D3WaX5deREvg7pGFuDq3qO1J
pGx2GrYShglpsx+HuOOwN3VIPZyTYv19N7AjNTS6jLS5xV9zvdEMFIjlz5l93KjF
+QAVFjP8vvRrFsplnoMLZTaCA58MXTrhXVe4OqoXz5tyWq2gRGmVCsEHrXpvT7HQ
O18p8kBZP3I2OE0TwayJQzegIQiohA8vMIGb3c6tJjEGz9xvAGCAgi4zy2ywnTa4
MYlpOqGyoNeomLGwz+oGLUgp93mIPCdBouyJBKTJaLg9364UfgtyWzSaaC9UEhF8
LbqPU7X5RQulx1409wl0KtrzPuCsax63fVsZpYrdaRHIGp7D9ysEBwluTfcb5sPA
LZhnGeJ9xyJjlAfBekvG5o2mceRGbbKr2JUMVa1Bt29hJRnTnDnjX1yPKez90cOP
PXUbhBC5eTEe683PRG+uI2qNcJmuBie0hzIZdHpl3HBnDfvfOx8nt+ktlkVNiDZy
c8mmMeCwWPMbxX+9E0LbUz+k1XK37opPIphXfPHnFclV4Qz394ELpaD5R+6fqans
Gqt10W/NwU9OZB628LY5iheNU7XXwOO0+jgZLF2UGp+xalnPX5LzVPtAeauMOrEF
XHHKNOa0BoMsUUSdyRMcjblU/M49rTo7+64QSopffxuFAGBFkk2HCZ3/39XNSIoq
uGpnLOZ57AFqknSh0OJogxqnCY1XHxiAkO3redCyeHXrJq4o7dUHs09JFzx5nqWC
uXTDNtS3XAf6dLH+Hoozt/DTz6c9M9uLXc1fzO5QybI4ubr+o4tMUN2X/GLAslHE
wVeFjcLbxSTTFiwHHrWhf7q00dvnTQzwM0TTq5plIiwshBhLjZcsHC4PnW+QDzVM
PXyUPIYbdVwwnBPCp4MR7biBYI4VJY96kjd/vgwq/igjjJkHTjpAUAjlX2bh3DFs
mXKZESzCuPRd4PFObOdls5Msp2n+7je9Sls/hNmNvF037JbjkRRB/iWgvAw5csAZ
+7xa0Y9oTGGDb6Sxolcafb/RNQwb7xHrfEV6+bfLiTFmCaq0Twvu/bvM8g55j3L/
rcdBoXao51aZD2w/3rAd6DCeO/oVENr60EL68cLQETy/DyMNCEx+jTMOjl+zmoEH
5QL4JincevMa1qqyc8B8DY882Dl1C/WI5hKRaI7q9XwB0+x20EaKtphXfuLUSQPw
UkRIPfcr7PCTw8jj+KPe02zyuPgfHznlPYXd7LvYe/XEdzw5GsNE9EJlApyyBE6v
qlz+5T1oy0D+2jV+n6U2krIOhoKC7A+nU3qm+3jyU/1NFkzt0+njBvjjc0cIfSXE
RNueug0A0Jtskg9FbWZc2GEVlSueZa3oEWnbxK7G4FsnhrcRHeCwqx9NYcpE6fXC
lyqxt3J4NayyNyC4FbEizmuICMeG1+k3HvTBLRgAa+Zca4RslSF+wnonmqkIKL0N
qqjJ+fAhQ3GFjfyfvthJl1rvxGkZHRM09vB476OxnJ9Dr4oECyVAkzu7DrQCqDjz
Mb7LRxL3cX3/gOOC/gQGQuKRWzbE6H27gMTb0OWRmOiddHA7WDafjBPk/4H4ZR4y
1YD/3pvJ4xL8lN3Epeq4vXx3AiRSEaV9G4xXCIDtBQjSqU97dL/dyUj/jrw2s1fK
wFBjmKkSMR6prkqIfsk3DB/HQITJts1lAgpiaXsskvbAWKNYVFllf0KYNv0iN3Tk
W9v4OyqYiebETo8UeD+QwpBfVffsNqYVgJWpZGaCAglvcw2VbZaiaRsZ2xr3y0E0
LkGGtaX0C7gN4x0CdneTSftPLJgdWseJxPxnJ5QxTbL6zKDkCxA7zJzJJArafBt6
nd5QK0gDphtbRwdieiXBcEOjThxCDoceewT4B2TmPvWtEs6YsixfpvwwegGKl4Qz
/AoqHDUIaw5wyEMaF3pgdh9KAl6DxywQauyYpe+jmF5KdYNkb9B/zBXSZaj1JOpA
ogWn4tJas7BXjTPys4QJZu65GtCMBNKiRu+HkwJoTzUD3W/tCR4RLhrueIQP0xXR
rSlg/uz7CS7lQ9UWT94pTIbU6DAWk6CY/rMwV79A0l/ZhUd5wlQ9hu2T73l+s7mV
P0LSiuJexNSc4VamU6XjumGHB99dYErc6xhqNiDF3jO5buWPNGzZmnqVcKAv1znm
TOh5ahJEL5trEsafWfCxjpXvUsV1UtpGA/IZUqgQro60tctaSQAXHZYJpDp6VqIy
j0VEdWOm1S+Gq8nwkRa0N+3ynbP7f3JuTIJM2O7NJR+xh65xSg6sO1uBhYNju0VJ
WdSvpq2nQjypKiP0UCWjgMfLZdmKyIu+j9ez66yR6niV2e8+QFfXX591bU9feRJv
b13mhcsGSBAhn6YwCHoWTZ/irlgp75Ed1Vpb0H+Fco2dEa0b+lyutU9PKer7SJd1
7EZeoM7bjcvkAJuDvRqSmhfzVpXqQLvWwqukAB48J///BDtQj5g91FKj2vf2ZvUb
DSd27hflJEqRBWC/ZRzYYKmdnBp4f48Rjb7Axue0WXVXnCkU5iLnlnMeQsBlxw3u
oI+cQ8ivZduVsQXTvjF1PE5IV8c31jV16DVL4uweV9AjJ1dbhZfZ4bvqJLGU9R6u
98L1w3WIm8GUF9I3t96d2YzMXh4MiZdbjzx8XgK8EZhM/YdpuD/OYuenXzbVTqTD
iuBfwlMfeUMxLyKPsk51DBKPqqA10Sz3CDkaOxT03wbTh7l86knlF80HQklr6eNz
WPNDwQpOxJ1kd5wGdt0Yts1rl/3o+v30AeLUzyByRExxUOn6Ywsw4X48Vjefpxkp
yMFbVuB9ofV0nH3HhFM7ErZfJHcZTr7o5WJ55iCbYNEeULR424do4oOchdg0Xe2V
h4h4ZoUVXGW6TC8dyE3ZgXXA1OOrSf4JvdIWhyaYssSV2hNmfmcYvCf0gnOJn+es
uv3f5V02GpYfkxQzsRdjBDnnPPifOt96lDwk2bt1eb1yhQyQyjFFYUWmcxMIaa7l
DxJKvtgcNL5cIe+EZbj5vGC8Xti16m58hCAncikGrKSG0i+GHxFDT/bzqo+tVoB3
/ORxgVfZOc1qwyAGjBTWJF6KPldh9I2/upsydZzSaXZJ3BBbOItAOru9JlaR0+RG
hvhW1qAnS4LYINOkFGQP9C2tX5uHCGQJTfeZpPoU9bV50u6UvX6nSM9gBKvkOmJy
d5OqYmlij5b9wljL+xgsR6TyENL5GER3LHv5f/QsISPElT5NzIM+blQuUVkVRnRs
3CC6xYLhCfhBbOxKW/65s8LqFL/sk0v4IIKD+Nxzudb/fVqrilrmHY2QAPhj6zyY
7d9H37Reo/DnEGOKOd9122m7VVC+QhwMZGceLdaAwTOCVygo90eqvPNq7RJ4YU6D
I9UEEF1NQGlsrhyCo0BT0oe2kx5j2kbosvUQ9LcJm1qf3ohmKDoska2Took3k1c7
YiyaaClcAkqlu+4Na6n8HsIOxQLz5vn5rHxGUb5CB1XhUlj+YhVJTWLpAc9PMzci
VCmJoxJmCc0lG5cpDzuZhbwB6H14rjPRlDVhyWMdiTelhtHS/hAUabmZSW+EmXI5
X5Csp585s4BqIDfNH5bBU9W41mYAM767D2ymfR0+jG0bqIJARIOt4yIMVkN4po6P
sKgU7REsCCE8zI2QECynG5lrncs0koPbe+BhppwR90RI9eZiLEb6ZGGIfPLPofPZ
d82nj/1viDFDwbfKpu/kgs5exBAF8IWfq6oa5N4KpU8y2u6XI/Iiu/hGIs0b4VIx
FtkseGgeLJcPJb+lZyuqURM7X8AM3RM4W2f7RUsX0G+QvX1wns9UdmQ9rbKuYVxR
Q8iAWqQ11xmeGXmlxOXHkrNpqE9zSvYmEDDaLlN3ikL3vGGkeTyHILhjd/LZWucN
nPgm3fTITnlwjQZIqN3A4kuXEl3LsnZBCFaquLE8qdsai8zwl7uF7IR5wxyVL1Iz
lBQ/OWj2SMZ3r87EDjw3GnB22i2vaHlRf6fCgXbcmcbB2mgiJwtSXkHwp1gEn0ot
kRexP5zsxHHNbJ/ALhi0Ils5bQY4fGuIUKGpDLso+rxzozySzok6NERgIOB6w9L/
eakLjTG+e8mDfuT/qhNTrwRdPRSN896x60iT9t+LzSfRQ7YahMemWe85Q431tefy
+o/cUibFREVhrS2zZnlnMwsBB5SEDJyqShuSnAnWYboT+oIQRDyiYgcOb82clHsJ
GATd5JVIiVJt3Oin3IIjODyS+QGS9kJ5/kj9l/mqzC0ih8eaUuUrPI+1u9zqIfYI
LmTZFIRSpFr/v+m/T1AzC82gK20ZPMaLvYrK3f6riSYuXL5ns8dPtzot4/IHKi4D
7/spaPCxaY2jwLPM1trVUJKPeWuJINlR4LyCat9afSgvMlOfkwBdos+izzVFX9+U
H5ajaL0S9ILuRLgg+gqpIzOULvXE84kazIy4J2cjysqO4KvBmi+9kktUm1CnFFvI
6K8ECp2fuSp4Qo9EgIqgTHH1RNDOi4gVaif3MjlpdgnUtoX2nSwctAwh+IhmEhac
dpRIcAdIZEVSuhXuWS8ixn8r/VJJ8SjAtXNhyFwiiFxupHBYG3yNwjootyI3IRvS
S03oOTUfpeJFG2IR23tjmElHtgd8O7TDunggnqBSHograJkgRVH25jA/5uOrgera
N78oQDUcP15g0Xakci8FhpmjrspR7MyZHRWjyxteWBvVLJf9OBpcYfy7ChVwflRj
EhdkXIxkafhbafMWivWhZQXIW18IxbiM5xemTd8WcPf3XTFqhPSCXw9Do9ID8bWN
Z4+BE8zVJ1n4qgb/MM831DyxFGgtgIJHaP53qJL40aVmsOYdxyQ79seEBfDyUWHL
500qiW78A0KXTg8KZODF3X9S4YViCjc67hlJZJWDaIi8FUY2kqeoqSEC3IPxHhtO
yW7cpLaQoUtPj+OmquxjOwup5M0jafcbVt9vFZ8JyUfC3e4hhEZAlpyfJ/mGaqnD
92EgaYWwBQf/St2dopsEuJ/xmj+9JJppF0eeGADDlJfyTnLtSvRDQueSOTu06LwN
sVbVo4Zy6VKgBUqjemmJ4L+lYhKsjppJZh39QCBpX7bo0C3OJAkIl8rIh3NyyGlH
yZfXHOeMdD6E0m9vxos9XH4LieVZfnJjdSKzHfgk3RRkh3dJhKbrYDZhEW2Giz7A
7C28sbpChLeopLmCGlP0ggzmVkHz2IHqCBz5atU4OALAWaeYXaA9fT6cOGRcihDc
scZ7bceeo2vuaI9fS8R1Rs13Wt+y0nNWL/n5IxZQNlOds/Ua4TtXsojB7TmNrz0F
VUnSQ7oo/TuV1vChjO+74PUWk4qXfhTiiTyzokpd/ZkIAw/kd5syBKgEyJYmy6zP
qw1PaP/kb1D4Dj8Wy6arhYK8P7vGGEUG2iLmSLCipgcxd7eNekXzuu/vy6dudD0x
O10qKDnvqc4p7NF817uQl2SCNMhLETWy353b7Ho1BVkNGp6ZcTrsKfO9EQpnX4yq
vPUvLXIOp1miqY3owfElXXMsCzw3GdfZ+4iR7Cv8T0wWIqIR5m5OOCvlvBV79mdi
pwp+xMoqN4eE+5lvLYQXDdcyHCniMD6Xjw+mQnCWOg4JxigXgxdVb1TecuEW5cJk
nGZi1IPnW2Xw4a4cprXBfBv92atpLhPWPG7IpmEGqD096QSWm4R9BAFasQ8Tl1lh
SwK6ayOAlSO/sKMm0Q5tugkt9jbp14v8Jgr9SzyDq5X/uaW5Lu0AzdcJ6zvzOg5G
9o/ymh+HWzTnZYHuq48QnGdKC4Nmv871GCaFgGjg1p68zAoBLrGVuw6Hctct/lxw
F/X4SoTYlhjzGoNgShHYv9EPT/CQxhLU7Xctrbu0uJ5eBopvn2hWDnFtdl8zRaef
0lO7+8lbGHfQhS12UGHBOCbg4aixUwCDC3u75lDtzMEavR0jFi96s95MfGIhN90A
2dU1OwJegrWLQKZKUPoxVBVeKyHopMQMwHCNkzenJNk6K1aWuOriTDPjl8nU+jnq
OAerOBhh7fjyVAN5pe7wnBOzaX3bKex+E6WAZwXbQzwCZEvqPWaxdepQoof6ZVbQ
I3ECfkfYdAU5c3WpvOnPp8YRmwkdblPhrttoQOrI1PLFqjirJvv3/M6sTkk6UTSP
Xs64WXppaG84OBruqh3h9YKQIDf+ff5HneQ50HYVlf4/6hxallJ7/qwInHAMaI7E
i04LLXVzq6Cuzcu6pcdNhLt15qTAd+g2+Y/JsfS3iM2dkTMgtqUdZWK9kcl7cyXQ
BpEVolBZ8BMdS3+7BKWtGYBSNQ8Z/3aBJ+a+ni+SbJ0HRbm1VhZlHSIArUVUdOQV
9ScVoHS5KdNmZNyL2KwUqpeaS4t9O2wSdeurBt18HIUTgRZMcceiDstwaJykO91z
/iVtkVNpBFRT5wDlRT+iCJT6KEas2jA9XFvzBaGoRN4JUz4qYhGy4GQVJSVwWX40
TbAXvFza6b5UZbyATTePxD2UtrwymozzRlr5D5k6cWyAyslF/17FxFJNx9lZLo6R
J8if+6Fz49rpnwZciaCxy7X+pKpJ/Q9nfYPBwGho1A2i+WJEa19jDiGee3by/x6K
xtTqZ/a1LACWh4HuapAmHF/6SytKAst5QCHvabbAXdCxjScZ1sz1cWh18V/+0Y7Y
xurCW/YDkk1yqU4NxX1Dmc77YVpIR79GooxD8RJaaOaRBAWr70h8d4snvR1aophM
2jUgO9KeR9qfJoYv/qQnFnEnaAKyBNrCmW8Y5C/M6TJY9yc4IemzXezr0GfT0l5m
AowowsO1bdzjhz/fuIunmZ1qaydqMqDFOIXsghFSSgOGORe8+ZejkVRBaEVHyU66
AzYvjm1SLuMiCAZ6CdANeNXSfw22oho4MI9wiNHTnGsVsOXDTRcLdwTCkx4NzJaI
ZiewLRSTPO8eOs5nZDOqwlO5/7PIqmaQk3QJv0MykdanULDEsbQKXktlXBYwO136
I8CqdcBYL6g3kws3PV8MAlSLz8MtgjcCg23TY6EZAq8asUCCh7V8A4wdxy8UnpQ2
R1wtp+QJjTnJ+q9tECJX6wDoKVMW8g7CyTkhKxhN00qba4YduQP/CwndgCSATXs+
Fo+WObIAUxiKHZBdS2zp2yBfGN0z0ED2AT1SdxH1pmrwBBPQn4TxgX9i+PrHX4Il
eZCMNM+4n907pZk1bOuxluI5MKyyrRzUxEZamILfKg1f3GdMCI9FHFoyUG7UA8fw
8cvuUyBoeO8C3akYp3j4CX0QW8Nt9b7YQz+sw5dtJUVHhIqFi/rqLkdmaedacpT+
geTsmVgYZmlhal6F6gSJlRPpmlHEpiXf6THkw2iM5fjjDNlwzvcN2fvs7MLnQ9jz
h/BWSHfgBMfmXWsPQlVVbvb1MWlLDhPsuwmsC533K1ysEHHgI+bziafWM/ILEnfj
q7qgw+UyXIGKvQRUaPi+jNJIRxGcnJs2evp1mq96DrtfiJf4ZCOvsFiyklxXFxYB
+B6lSBAZX6FhFdrtUmQ/S5Mu8XX5HuPpXT8JT5Y1p/ILMnvWmT0n+KKcqzwhfYhT
6HXHArmzvu7/FFur7mURH0vbfYZxjTRB84zioeHkaw0KTSQkgagrOpfThigRicTn
KWJkCZLHH1akEPA9PuHFzSiQ3nMDalYo6jEGHb6KM0GSqwOxBuAoMRPn4VuMB80r
wbdt9DMQ7/vOLN/VX3uPnwh5x40G0r2YIKvJkaj/qMDZzrA0rioOXkhQNchHxOmJ
wu4Pa5jtIhTEO9Kdf7bCSRy1cF7hf+GdHosSAp9664QtT1FjIsQW8F8+FAQ+56gY
66Iv99y2OP/C8gLKsS99mmmnYf4q7x5vNKrCZqsRMTKpIvc7iPUJoHRwy5XLI1NI
ktU0+tZKRE/pQLKyWEjG227kv4rUigQTW9ni/d0KWt/vdz0to4xDOdXyqObM+k9W
vw7QEpZMcur0Jm2ytTzZJkxHipmUcYnkQ2dD9p/F7x2oloveTGrc63va9xfgjN38
f5ULn7OYGCx7Fy+MsQ6hAaGDChPgu/d9GbYXitnRtMOzCIx1iIK0BVgJxBfFeDeR
YcrBcK1dupEzOBacdwJecYlhL+5D51U2E3KK5iTlaAqJB9+pitzCTjYpzpnr8cg6
ADX9OCNKc9yi0wVXJ1RCIPPK6NVlcBkLJKgWBpRFQj9lC+jtthC6mev3lbctfyQl
u1NG77+FTQ2pmuBG6MNDvquy8XCiprB+vXHiZey2+gYPb2Weee9K1RwBcSqGsKu8
yQ9PUHyhSE9RZZgY9HIREIY+QLcEJd4rfGse/ahRkFVtztufaMjs942WV7fNTTKG
kzMtByib5/L59spHrO9dV2OIP1QW0DL55sSo2IfztzDENn1oGqlvCpFgUh2fvaVO
quiwOMXCh3WB1ZakSPKNDhqU8Sicr0I2QZUko5eQBAxh33xcdtjfxlVhe8c+iqEC
EyrJ3yTA40dvMgZadiV/wvC1HsYbL7iyELMa8fHaMDSRoUW/bwvpYYHOrrjv5IH3
ApYwncHB43GN2/vPy/2gCY9qsO3t9OoMDRYq/iepoAoFLL3HVT89sxksAYbPB7jk
Zc8dIVpY3H5mNY8fscYgVQacwHus8/CKcGjnrhUK++ZKVCYabFDwBc8gKVowFxGv
Fo6wmuGaqYeJM9cXD7hIrvHaobTSUuHEsOLuwX01gQeG/nbpOe8mE65UfFLI6ZWr
DMQi9AlcUFsqPgwwUYyW8acf5B4x+RrboxTEhMJ9j5TVTgdUdc+wYZ14zKYz51Qr
xHy9MWucBvbq/jxyzt4DDUEsUEO0fUkeAZ9JJQi+zVAg/22ffvUO+6YkELqs2n9B
HkKLuRGBd5hZTZo2MEoYNLszqKXUQ05bmVZ/CLk8T/8KsIM7fIu0luu1E+kMZrIH
acDMfx87V0vAk3xQBKrDlnynxlyLL7FbOAH4sjkoGY7HHUp4vu+WxsylQ5mLe/3J
6QrQfWyQBN2/qZYPBXUlffnniIs7lO5EHZl6Fp99TiJda/8q/g0aACmrlwTdwpXI
hNwunKTwsHssEzDToOnpKmiVe7xjDkG2TjQVDzm8yBPMA6jpk28ITG8YxpoFN5Ww
HB4yAlVuSNBbFVi83OwZZGRjyTGLdZ7ucAbnmB9s0ktaSKb7bj5mgElkpAhzowui
c1TJ+/eGe1OdZep7txaEcauu5XI2dRjZ6BoZXDqNbkD+Px75vSZFBE2jgBj+VTJ9
7+X0yFLLm5aFJ1z4jZIzXnFZaeJDg8fpoD2kX1H1necND8q+FBy4jhv7RBlIdMpa
TxYdsJgxz1ZM4QjBdGKmNgfvsftgNuIW6HoSxZDaW7YHR7WCVNlmS6fVkQtW8aGh
UtrMTzDcsIwP1kSQd2Exk9MHkso4b72hUX194P8ItzaOFd6BYj/eAYNgg6giIxKI
Vj7dhu+mLPxE1dvYyrll+g==
`pragma protect end_protected

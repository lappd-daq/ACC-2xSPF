// Copyright (C) 2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std
// ALTERA_TIMESTAMP:Thu Sep 13 06:36:53 PDT 2018
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Yyx5Z6E4Xs0wUtW6rzEoEx7Zalmf7j7vY9GpTUoHtYkjzWQtJ0izZqjphEPuVNBO
cnefPXLmz1usJq7N1nNa/2MRUJLlub55T/sV1N9tNV9yYztoVrxZeY5/7OLnxYHQ
h6BR6DYTAiTLMJZ4nAEvi0a5nSCX+QI9d9K5XCfbkgA=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 25648)
blPA4hEEcaGNDp0NdROaNP9JY46o3nULUOnqzDnVIuH7rvdrAeZni8NXrl8QMN2C
Il6046NhAl1kDZJFgJO6kGh/mGvCPLhZz9LMFtHcKcKj0zL1gN3aZkcjkwSLY7Up
n2y6Qu9AgyhfLyOGA+HmlyODQtscerH3c3qPvwn1DNcS2nPdGT+3+5du934pvbta
RTQi4orlOJ3bHPz5kluYSSOyOmKqKf3CUC7jYD2sbULMdzGk0kdRGW75volPcMJD
Jz+k3xXhSAM/g6K7Zqm/deJDb/GtBFQF4/iCDsOn8+6Km3fG78KrbAqr5ETlHamE
9fTQeUpZQETe4UCHWH5SVPOXJMcqu31oYs/D81gS7p8j98lj3oOTd1onZ92ou8tw
MjUct12gvh2Q3N8ZpLxeOw6kzzoqt/owMNYT13tfKa8uNepc0PKQkazi3lNtpfka
5MInXWC2l2bi8nMACn4gLAlMDi0XuXKfdGHSnOgJly6+UEdlIbc+Q6Hv7eQDIGMY
AwlwA7qQtjoUoPXah7y6zTq2V2HFTEC3i4K9XhRXPAPcT0n5XK3eI0vHOHRkxF/k
LewFaV1nv/k045zHDBFVN0F5a37tp+Q1G2k8sEm2UcRBEYG4gmjrLyfV+OGfIonW
iviDN7Hij20r3xj6aSKGNtdoQk/rvj4wBSqJGWg4VAr65cdYdLCeZ7xrd2m6j2/e
Fn6aaGMh0C8r16uggjUMC9pzCNYPR6S3V6ybvFbTPzTZkobcCa70LHl3j6dgrDLs
hSNybu58fAdycobb2C1TnexSWTQnLbEhUbAAwZFTNX2x3Ctq+KWsag7NBFy8W7NG
tvRG3pahOsOSDatluKnj0L05VoWHZNe0HddkjT1FA2Hyuck9eiBt6NU2ogIR7XnR
6rJe13sKfmCr7d5Q/gclc6deAg5fTMUlNB7KHy0m/nPkL/UFJwHMksR9EUqYhvg1
T/6uGIMRUVrrdInNX3s4Nek0cen1TDhZlV61SybxU4JsInvHq1zRYTRpGr5m9rkb
rbjwi0oJis0KOxn0j7vT9UTXk20U8CVF4/APetyGG3j3lBcwuUiTIUFrAojaSFjp
oV2GC5ZCbpfwCNJkW1nyHMAceNq1bnW7SEIUWTENPz/DT/5KFnsd4buTM8lJFxwR
NuNwOhvJuGg6PXOf+Ppfiq+3bgH1FDFZMmcr4bKUtR7DS6CJtzLYrwvWLoidStGO
4zQGCx3M91xYNgNrCUkWHHmDL2mRxGz0nin96qJd8ELEErDSMEDqetB2K9xRE7fo
I2noZQupljZ4jw7eUChlL0XwPGc8eytAPDDYcFD3FDgtjQMJVfIUn13ZbwdQVU0Y
2obSJHHAp35SLjps52vhD9+otCrgFfm8S6FszvDNGQpf1Cz+dDqCAP+d4Y3ZOzmY
xU1yRaxC1TqSPZP279dqy+OLbkBmTH+2Mg8NzuebRu7JueQSWieFuvX7FJGgkNjI
lGzDAkw+40ltWqPDglRrC6DdCVe3WP5n2Oa6zR8bMkbS94Ho5Uus+cqMWUfj81BF
eCt8SP+kKuGhkE/j4evPbZI4xbbK5LolqxFl18O+k0Lgpkz6FHdm/9E1+LWb3myH
qj3dgmlk6PKnSZ5YoK0FAnx+FFpCTq6MiYSp+jTmLswEYwn3VA0sBfCFd+F81L9g
99U6ehDneHo3HIFkSVSBoXDwj3TpUgXF9fRHrjz9d/GKFLCUHXjM0yz5umiPR/gJ
XrJRRH10DBhTpvgxjjVg17eOihegyZ42vUHnKQPelR1Q9/6oc3/WjoTi7D6q5jZ1
WgWCgWRblntMeLItS8F3F6tKO61Z18nNun0IS4aCGWEYlhmqb9Oe+4Mj5NW71Xx/
ZF1uMs/73C8lk5mVlVwCLsHzWnQYhv4g9k07OghSoQH+PJbFzYS6tKpSGuJsiJYY
Z2NFi0k7si8OZKNpJ0PwZM2JInCQ4AKjNZ/blyalfH1/pSZLtcYNS6Nt0Sv5/fLg
GYVOpQZgVllyPgOFIU+FdIEw/amCCg3yKbEzpyCqNQyyFtxsdDbW7ReNapcl20/1
0N8CZr46Mh8vcjZxvOTxeIF4dkMHGQHKF0GQF6WEKmyCmhFKVDuVtKJznBlhRZ9q
5dVIGi0y0spQDx9PkqjUkpP0KVCLerIgI9/lOrRF3api+i8bMu3fbDIezPlQaPrQ
TInG9hNsaEM+B7stePpCbA4OVpfdWPfqkotrdwo6zlKRE3aMbuk9l20OuTj4tbts
QvEsnjYE2E5WqI79NHnOyH22SpwzEF8kqCf7EKHzBXjmEG/OoH+MzgNgAGJ3/I/W
T+UKSWhGS+Z0yTtl2KuLeXQPLxsmEhjPXwm6/ktdUh2MUj7GOyPKhYh/RfHdqAK/
syObVG93XqEHn0JQkX5J/fnNIE3KW3n1q/1W9I5OCHI57xaFWxL4378WmzL2eKQd
DMBjvq0gVIzoQg6UlH8vyMkZYd0ZpLXM97U1Za7jVDY3d3ICqlLESUDXn4HvuMR7
nQ2VhR7DN5D/2wDHx1d0jxGn666l8q+ESSA0s47WNTKzX+W37PETVjpbBedaVTET
tttOegKZiVjVWo4cl6xwriPD71T+jWV2OuOx998p60sZ6Bgc6YlLWT3lJmbSfTY8
IODNFc4CFn1wIZNDNiNoUurNdX9gyPNlgy8Kj7fioN9baqCSb/rv+J3zOSazjmXr
ok89J0ipNtnZ9r4kzmKWmgOVoWWulSyvfBPiwlyHoez7+PUBO/qfH4rAbZsJJRct
uxwAXgHELdoHjUTRV4SZjbWJRZfmfYpgtUwa9GTeKmtdMhy/BGqpQ7RfcgOQOi2k
XtAjBo9TaHfyh9t+7M9bIYIdT4g75x0SbVC5BXE9bzkS1hNjTBcF2J2uQAGyKR2G
FEan5yLnEvgXkh05MlleznsXUi6tDmq1dhztap1NGjKb1dXzVRPJWbJrDMztbKtG
apJPub+9a4XG/zEha7dZA+1K1YBc1JfwBo+KsGg4239CE8SdN0L7pdpFzZtRLNPN
dG+LLNaSdFYqdY52oZ37/50MsoQ3ow0YiqykwfsBihJDoUeDIl6Wr/mlHzLyuQPM
HSBObyc78ks3n7PEuWLceULg+wz7HxK2sYwwhA6twLncw1jmFc/kv5aRU5Az+s0S
iMogCBBsobM4tuOUfsBtcvSBuBgWrepE+7LY6daSvv5shYpVZNC/j0232npTH7HP
MQ0vTOU1q3DkmlsaDyigzj8clWl+qz1o0exVrNBoyk5SUV/rusSzogTmdh7H7MjN
wJLd2NFrVxwQBp26+Yfs0Fym6V2SyPB3tvj8vyY+rbf0ZdVhyuxCnY1tj/zAsT69
N/uKGL4dLoz+Yj7+Nc71ti3PX9FkoCQ8bmBOQB5RK4hxEultJvfCsFoY49OftFqj
vS/SfDSe4P5USrcCzxqDNutEi3bjrZ8rxiTGnahDarWgZF6aAaU92a1ILA2ZRDRU
bpsmC1a33j25CLUgkWrQDzzsID0QUOPw0K22gOnRvJIfTAhwIh+IYSVHXeCHeTkN
iLOGLf7h13jEi2ROsRkHCyYtTGQbEYGuQQRd/XU8WmoVtqqP+6jNqjrx+NGc51qC
PdzjtAFyZHhnPFcIKx6i5XISqtnZn0khOGQJnUgenCkHYPsbYXHja6IeQR7DIet+
09G92rn8dz07e/aQ4GkKb16DAr3PlBS3KKV3UXX1jjUVqlOgzlzMSlie0aVgJ09M
eWGy9aNM64G5wXe6fokHDJ61+ILdipZQ02uoaGut29Wa3NdpkHJFXwLgyZL8Hfs1
TDoqfrshneLTgiRSfEUf3jUfrqE8Cl9brk4bahgfDSL4wZtAm8WXSvvduobwpwbG
nsKO8HwDMCnzZwT+9+M+qQjtLcjvOzBU/sF6P345OJOecAVSc83CTzOwv8SmgKQd
oWkFeDSsZK3kwhEtCORDAJrZ4INjq+F7OwF1bppp0bie1i97dJMPsDkibxGM7hLs
+z1tk+g3pCOZGrI+xtrENLQIQHtHi2CVxklz4buWXcvRLwCYil0IbeFc+C1vuQ+P
gepKHmj6I1Rp19sPTS7TXXInbOYpS4gx3p6v1rYuMdFMFuWyozI+uJR3AZQYAbiE
0niGyOKZ+Ji9TtXlR7MuNjTGtfbXgnvnUBkp9mocynkHXIvYTw5XfuH2WR3ZiGDH
opASoTQgg26SADLCcSD/BLmHW4578HWbHQh4VJQxOLlwcs9nCDaaflKLJzudIzAV
mPzvHyzjqINltw3lJNYwtjWKW79TlWF0/45nGxCtYeXlPPwW5GflwjYlXKNMSymv
6sO+GGLUFJauPQe4qNfr//up+Fa3jzP3mr9sECfZPTAKy7GLhZsN3SJMMPO+q0dp
MH/YuZDjTRbkyXcQuIwiDkjErh9LEzuJfWu7QbipG5xoIqIWWRmiGIrIsxZj0LPI
C67XE/93lztpJhV6iBzzK1o6NsnvfoFFQK8vGa7PByfEU56lQrhDwZxQFU9EsUct
5EGUMvnynQzxDPlCKB0eu9kb1kS6w01MyU9OEmOCiOCBj871UPVslVBi7MLwTZjD
6tyg/W4JRvCg33Vc/ita1GPPNiOcXjg+eTDVBV7vgxS1V0Etk4Lu1A/Fmqoxl1LZ
zyUvFfrv5NEdLXu26UaEVZC3lpfcGxbIg+dkhx26MH7aq6/qHduQupANjG4llpYH
PXKT2A4aVQvX5gvumz/RvauPEm1VqeSqVwjzff+orqkLALhzQtTuPrQTPwDqGnFy
2fzad1r0cA5Hx6Nz3Xv7UxDpvg5/d7jgWiwqHuaSKxRUtXvuznhSST1OZO6Bui12
8yfiTAjVOfQXohOmLZvO7H9RHVJ/k+2qKL7bKS6OD96NGSiWa2gXcaf+fUm4j92s
JKUssaKPY5TgIB8ehZcdtuZMmxx5iQJkU/IRJaMafFMRpoEvw79njNEKpF7/FI3A
2IF+qxm1tDJKXF+tjnq6VdY+pOrM50tDhR+JBsScq2f3RaUdfLza+7Um4zJtjKuP
BnjcUyT6SrMzLqkk0mML84OVBaJ1pJ54FYrOG+GPlghggYslhbyfCt/mB0zFwhtu
Oz6QCi6Kl/RU9OILqsopj9koeYugXr/SMXiesOoCffwTh8uCeyRNfHxaIwFa+Q/E
4a5Y2a30Aqznpyf8ETFzSMMiyteNVNdV+68Ysyq6nXYSGsRPNql1zfQVqPDni8tu
cfPgcdh50/cuwxqcYnJP/pTX9NxdDX8N0A5AGc8muJLkBmYhk3c+DJH1ZCRITIah
/J05BrxZcol/BHPQ1hJMdVPg7tX4qpDlOX/A0hbM+3nGaj7tVHW7dBH301nJgtcW
xr7oSlX4ai7JYeRBG2j6gN4beSurkDTu3H20P65yHkSW3UobnvjHzC8u+f6poZnn
Sxr59vH9SM+aBQyfNX7vOIC7IoSnA4ta58Gko2Bk8yhDdyfSor38GoRe1iLuc3gY
J7cyr7bTs13DX8U0Mlfb8zeMjAtGz9O+TO/ttrWlIFmSuLc0It/8UwG8pgLhg8sd
AzcxwGiJICFU/ZnEKqwHymA5Im4MtvqYGYhNHV2Qt7OS68DEZan7zsN9Muk+hvBg
xVvGPbJ5mafiUzvpFegqdmf2q5GTjA/pLW7D/YuVAlSuwsjBXNSWe2qayDgl1NLG
ixFCsjj1oTNRnd1DkUjZpWOWYdgKsB2FPv22K72QhbUvCGheGFm0fbRzX2LyYwtl
deOjZ9acDKQeQaTKHZmJjamlx25C4inDxqwuh53/gExEJEoGk/CDFizBVnE/wCOs
Ga7dVEXNOHpu87mYw6FuqvRMAxHlJPwbb2QSRB1uBJr118wH2DPcy1d4Uuodyihw
XbMf9SBVftuZk1qyD6qDL1+aq7jlwQL13vmpXTzxITgBkAKQKHapzTpLClz9tV69
nfC+v87kvfuQi0cX/YajUdSIrhShED8VgDgqO7/n3GUeAL8ikTA2bJlU9JMrNUiC
teSwrA1Qrn7W1Q+f3XcWSvLlNU3fXjCEbxOMUL63ImFUEgTQ3QdMdZ1y7cr/M+2Y
Y5RqkcmwGod+Iti0nHQqcideeh5SxeJ0wl6i2G9TvGHJn2NJPgIeHqu3Zy+Rztty
0D9lC2z9XjTpJECwwAr2sTXiV7wTKacwbhzHSBVlH5ow06FzpKmW+yTOKalzR3fb
uT6Hz7oTsjlUdA+L6HuxK1f0lc6VYE2UOlcZuisdS/cHAYd82+KapzuduGyrvnqM
bc+2qlaR/qTJn9P9sfckl8qDOqzUCqJqIoch8G/4Npjt2jJQqq13VAM3lALdbibX
qrCdoY5vZnhBn+ckQz6fMilRoT/mZ+RkPviYN+oArSli8DdY5gI1/Sv7m7b6p4Bb
eqRztRolBEtbd5gf7lLyBUPzp/NmGBS1mLqz5og5+ZDeHMKO/qpecwCFR73W8RSr
W5Ivc1r/azg0W9UuMTM937eUiZPOG0CmeRpaogmflsn2Zv+adXtdmG6j97cDQHU/
3bJphLlpA85AMffC86znrTZN91GlBY3EiNbn7eVU7Aux9eC40lzwSOClL9LLnMt9
LZ4Kax23uWgGHhyrO36Ev42MYrNgH9itSLVyLGKNSztqpQ5CdRmCSmgaaOZZEwWH
wyB8FQgksmBay4lEdEcvINFOO/tYpr+PbaMjLQnbs1nJOfmk+evMybrz9ov8LHCp
/uXMc4m9D5BNRYd3wZTn4m46izfcYuzvIsCgpfpmhGKML2UTxoi7Wlot69Huulil
lcuB5/XGe8ooks+DeUHz92SzJN7YVmekzQ3VK2N0ew5jXNrIy9uAf/nlofRTFV8g
vBpf47ww1F1vgFtAGZ2Xg1Ak4GSiUJ6X0RfGC0n69O4n8raRLTTfqViOuGsb1F8D
KeZKtjqrzIboFN2ct0PgVg4W8QaJdPvkV1Tstr9NkXd5C27gLp8goqe6k09bl4zj
VnSZLB6wfXnikMBYH8sMBhlECDlRoga8KBn3M4Jstq2h1gg1DgyqcYVLC72mz97k
nhSenc+SfRrL9QsXewBt/TN83royaAu2JH/V45AKEZqUYwy/f8NaTsPxcHfnpQef
eDthcqTSGx/2DYw1X2LUIbbafNWAmoMYgSb224fFfK6dS4Mjf6gtlxUL9l07iUsx
9gbeCaJvKHy2DRQiwK/q07JWMWaaU516t7sKG/amQkzyVthlFpCf11Hk+/IX234r
nrLgj18JZspf4vpKPSQbGIYZRJAH+GFBJezIlqvOAF5R5qB+fMoDooBu3FXCzUh+
U+4i8OworYeuTAj7oZdqxKHWOmSzTYEVBJqqeAFSfRj/YvJ/oWKnP9a2Ul/9VLEA
L3yqY6GpZZtJE2iscN3BdaLWHIIPTSn5jR5LW0LV+V2YIp4vbPe/CeK74ZjtCExF
XC0fOkNeR5Npct7SMFQH11e162kOf7thVM/YV9OhpsU5cH//vNqD8Izsfnl19EH1
Xw/M3GTAXTOk1L4tqVhqqUMbn2l46tkVyyeATd7RtObkDce9oLjmApGSEu0u6YYG
nazJj3Ssf2B3cVWZKg6APA7HVbfG3Ywc8UNi6cVVr0WLxU+I+9bCIOMtQY2FfjAD
KqL+gg1I1heOx7R+FWsRif51psnZCOXnzelfgm6Aw1bVwd6hLM6dEpjfAEkaNLBS
99L0GK2MvLEWaIqAn/XmzCNj+08vJQUnXa+9WMv2INCSjUOLkL/2MiupXkTpYZ9R
4REhNzLZeYUGo2LgCqkWdOUSn7hnq4fOwLCuUQc0t+RCki5X2GG0G50eOo7HJ/GG
Gb7rsmFm3rxPH4+fcohBWtI0s+0MXWXIQfBAtc1LP6TUhXLpQON5F4K2JfZcVCqe
OeZxHs75cYY1RPui9352fNqpqWfl43Qh+xByNg/sZpp3rOGNZUM+xVNCh3InO9pu
geBlEeTZMEhu2GrGtN8n1jlcsqWqgUsMtJ7tZ8+w0FJXFPChL+CowKtTXdvK0vaG
5gXWvREEwEw43XBFYRguODGaLpulayCvkOFPELFehVIMjtSYF2s+rDttu3D1IP8z
LEqXtIcy7UZQF9E8xbYDhp9P8lT1JSaHTpLyF+i02PBytnVYwcjq+j9bHYY4AR+0
D5FFrulTRAZyT78CrB78Do/5Kkcj0gsnW9gHCHECb/yGXDnIMNFnDx/EVu457IMb
INxVJjhImOkXnlvSF5hoaXYVVt+b2zZWhy9GBFHI50+IEsRKY25yICm+30dTP0Ol
82ZrdlMn5aw1AQP2oEG5rzeLjtnxBmjIVh8uZeY652xJahyF527QpRJtDDJsw1r3
I3HK1OVL3CTyV0ZsYNBFzNAbKtA075DKq3Y36Gm8jVQcV38N5M9f6TCKFd3seQCI
PvuprevxeEphuV3GcWxR4+dPmqHiGAdTCGoHWabrQ9OmvVFJr05fbYMJibPRXkX5
qSP195P8+pD5Hq49ZnWWgAz7kwar+YBET8gXNE6yoSeb0Ak9t/0/YSlWFysEiUXo
x2VUgOcwsI6ccf1/h+sjavJyNpWF/v6zGg5t2oPOfmRGX2t2KukIXgp7Bu9XNLAf
C+fmgTnBKbWPhSJCDp62IPJ6uFFisrzQtTqXBF1+DBrP3CZOm0qHCaeDmcJNOeXB
oXtph7jDmMZxOLf1F5c4l4yjHGvLZ+mWtz3tnGyS0M319XD7criLZlRlcDgLqeZ5
VtMBGJAkjAcLmgPVOH32zTG3Trd71L5bTgYh6pp9Eiu3D2LxzBVmvs0U1iCicnkh
ezzfCpJccjv2L9VczlTeWlJ2RthIDDPXc2w5FjfW6O+4+XGcNYs7w9T3g5FcRAv9
EPjUkgDq8qP0uFph4EedOZwnvIjMkBWPz+lkLBfNqRTxE0TIu5QWa9TFLSbueJk4
sg+m0EgbZNUnBgX6agxFk6BFWIRrDN2NCU4q2B37kybGGhXs52ZOkJ5cDpbhfmqD
jQ+DO6Z3Pvvp9b02Q2z+O/T//PeM3XV5BzqvQTOQpRsHU9YTTDrG2FR11drsIs1D
6bXsvDtkBYSFCO4KGIffT8o7irB/SEbsppGFNLvTn6pBIgA5VMYrP+XFlt6YuS6y
HccZhD3KL+zqWo0KNdfq6Lw7fQKlF5FD70rrQhDJZIWbB37YdR74Q3siITkVLuRU
IaKlA0S76YRpDT/C25REVIpe3HW0Y/cxsYKHAZMW9ECN6kr5PJOIc0XHjoxKTj+d
4WR6CAbivCXa18Xu7vxSMbfNXymidXjVlQ3vIvom3MmzJLJU1HzOpD0SgqN7lbGC
LR9bv31OwlYD5Lm4sdpOCETsB3APqo3t76JcZoaMs0JQNxrIzOamZZV6ANUp+hJy
K6e/+PaURSEadWMZcImq28fQ8X+1D6hKc6bqx2cM5dNmfsgBO+eplwnZYoseqDBE
xf2Hmf0taqxnmBBbVN2h1sq9PH4zb/BZ3qE4sKSmXRDZ/qsXzUL4yfT4jd7jmcEL
6U0o3I+lrWdj4C+/Px/k5ZvJPujsWhWkuLmZsp/5CgC63Jm1wMzelsKd2QmjdilP
3zMiSbMhe6h+W+PvcAQzhI6zAEkGJF+G7yQK40VxvSYnxaIkS2saT3yUqDx9r//c
DCnTKzslXjrm+oPQt56z9qCGxrnnkr+/v0n+0TuUi1b67D6wV9FrU3aEIHcUcQjy
zJAwuiypBX2R7wHs55E8Xia/ezA1P6LZCkmR09gvUVfYvpXpXjMbeVvSgbA0RTWc
GazE6GkfzAMKHCreuz07474pCTpYvs2Y11AJ8oCEJKQgktzT639PyRPhV3BkT/YK
3qjUet3zYjAXLTAFbnSYaQMdlPUDdQG9CqOYjex7gD7wJjKB0HUALG1XMjGLjIif
t58pTUqjcmjheZCaCHWu4EzF+H/hzGJ+IGnqatvZJwBZsX9a18Gn9tEAAlE47fah
n95zAuWMjB/RS3O0qgtqVExM3KfV3JcFPzfall6sJwlM9qERUEMJSfOmVbD/mi+O
0npJHalb8Px5r7qqOFjZCrDK+sNeCg9kDlFqxi/mvPpIQKWJkCMJfXPTgQ+bIRYA
eO054hSs31GUvVWkBpgC7wd3+50awXxmitXMIYD0GnAuSOqOfRCqyWXNVcg+lJ6M
Br7OyaDBfNvoRIVqyNW5JFfr/mZJ6npeSRpo2908P+7sEnjQRI3abSx4XrdQRkFl
kbdZa8MYNGUFOs0bB8OIv25Hq9MzrS5c4DCHo7ADxvQOQW5Q4Z54zExROP41u2cQ
QzRFeM8PMW9qxRrVkPpqKMJlsuf2gcYIPqGaafGfhp3jQ8RjD46p+GyZRW5+nPvQ
SEvcJoNynrzI8u0UE4rkaF22t5PZB9PPx8+jic39rLy52dovoD181wwt+ADxnb/y
a4YGajZDc34Q8X4agpGgCHhepGjmR09PSt6cazoL1z2cHxM2oy8sGstcVMUD7SQ3
kDPm+rR4yoHEobkaPsRMXJhqbQvTVRprjmuGz3bNdWJhVjmjGYDDCraE23tbV6sa
He3SWrFWVusOTe9PtHQR+HEtYZfWtkWAFn822diGBalg2Dfk9O0KA1zEJ2Q9ATFS
vFiXxMlIbKcCZFxLCz9xGu2h2uC81Z/p74zdyN54RzH1a8IGdnBJys9drxAgeFwW
ySrKUHMWQDVoVe3440wBNQaB6SOlOSLQH1dSx/nVtWCVUFO2D1RAMwz/vmsE9CRI
6nmO9PqPJG7zo3oQKtEznt6Y2QD+DPqfoT6VcjzkS35wriwV4XTxp2zcjixoOIiu
v/qEUNAXbkFHKqPTwGq3CEj5H4SBs3APgVacpy9u9PCZRgA9pcO1RFYLodLe4N7p
45+2WKvnSndrVPnHjSWLJ2iRTiMAEEWq8L8jTJNbFNrTZVYvugqydDaeRX2s/tYE
ujJFXHMjfdQDTtePtEOjIbCz6MDMbdSYi9k2ELoPMiOqi24jfHKrAsh125eUvGqR
UKTLN7yuHP/ZvzRfUWUMETefPVj7M4yHhzj8wjS54cZh7h8kSNkoWpyxEQxUFphC
lX35MbCp5KOiuyRtkE1rXm7V9RxnGvZdfmSFoU1k2mdcL69Lfix3v+tiMWqXWz8y
7gEK2aeFzV03113JojgmKt1iT/+Ss1rp0GvcS+PI15XvJlEPtRT1x4267FMgB8O3
gtDVd93H3DHIs+MiH04e8q0t65u5OfAojEhLhjirMVFymwG7J22e5xi656FsIZQh
aFYawgrxVYCyLFiz9FSN00hqUOne1WkmQWWBXPLt063zzVXSsgTWm5+COwpaYyes
vH3P4ozF0TTCYxFgQSD92/ZSlzDsQAK89vKM6K+sJRHmcEp7ir9JZxO3Na7cqwZi
vQHzX2JAVIX+yioMBiy86yOqUW3eeZ5H8oygZr2WXTkd/m2bjv44Dm2dNqrmNkVr
QU31oJB38S2yoNbIYyY8AMSYle5k60JVlsI1wNd4Qp3VtNFCd7hUMZM7NcQOOmoe
3rjuZpghzrFlz7zvbfGLDfXcBSADUNGOcIzCRnXEMHAN9wHRF+trJOxrQdhFyrKT
4Ki3L4jzGdZHW6sUewg1nEvzA0//1CbgpjWDckmbk9JWZiL6F0P38gr39zPFU9FW
suMwtvcmkaCzS/FipmWK6EtcpRedSHHUeMCQyULWIYsYDiTN/r45uIvHHWzH5fog
QLwcuv2opM7L2idgWVc+KZ38pAHqSVQ4hz3Qkh3fb3f+bl1bs0CVEkMCLOHbiIaV
V8GldR27gjaJ99B95IrPTQ9i5KXY+22HzSxTHp19Ck+fyPqUoSVaqtOb/nquDOVr
+B5wbzF3uFPvAj+xzmAPccNNgRC6i/xxo9Sp4MyUbtRoAljzbkZeNTYuZR6Pvg17
EEs6baZi57xEi0nc4lMTHLUk8wuntoHegKPIglhiqnhtZx+3AnQVn2K2i2zg56TT
ZtMmyf4GLIAH2AitAn5GT0OQkoK1xBmYGJ+WIHwkZret4KCQdccTjmYEoy3bW9qd
ar7cif3d4BeS1GwqWJT88KCNOg4F/byWzqfCCsiDE3HdVWYHD2Kw+cTKYHE40NHR
wBlPjN3lMhbqVBjbXF5Q0rXO9xkPUfVYYGOi5XDXRGiUeiRykuD4JGDGVAFzQ1lP
UUt8vTd+AOJ3MUNxDjoyLubAb0TBy1IYHSxStBCRYn0N2trVLdB+eXprPjoeXNgf
sL1DdC4RLWevDr6xiYcDisgxdX/Hiv5BZdV318G6vHZpR6nT986e3AVup9rUwRwe
X2ZZNMjY2MUdn3NW7X2W3o6YqLjoGBJJxXuPtFQXsMDT8HZIWv1U6nYpWQtyi49K
BuK6bWmh26CBArfYoKV+9X6tMOShbdGY1dx5/Wc5agicVPz0Zwv7FMntSIji9xpL
6qoA9DBdigpxyPQWXLqa7YGNCqVaGRpye+yLmvJDtpRCc6b4cM5XvwPTymFGPSzL
ErS2Qk+rv/lle/H0fiC1BJZ7oT/BfXHf5RwtLsponzmXNFza3OzhCGxqFiC4Ek9l
GbbK+/IFTF0gxATCEFc2wdCGBC7DKCgUTkn00Wf0dXnMgQWC+3VALBahZUXLy1Mo
gjD3Jc3AzDUksp1rcbWV7zdXLhdx2emxYbkO46mHLj2we3PLqIw9PAvj5wJhytRb
qo4lFAWIX2nKwLvfOZw+0Mkv92JurKTnKqXnw2pmCQIu94S2cJQcLqBHL/awxUA3
hp0sJTDRGP7bdBMcwZbG5R21+clVk5IgrSrGMydzyJAaTede6yQG5wdLvPGM+QcX
G8wnGIklNcTkBl5EH4HRXEeF0k2JmZbT66PuGK0G+3Ob2fYb8KaFyja/nEq5o9On
2W9jlsb0Db7EyyYvjRbGIbGvkFgwG3qCl8AMXzaxzMMPNOyNR5zwCrFs4hRt2v60
alZKsoC88/wcEusLMs8t1mryWQyHHiF40eStcyQcjCCl6FqDAg6mTsMD72R/Y/AH
qob7uFol/m2YvOzEXKP38r8qiQCwBDMzETDfy2kSnVrgLrIhp5T3OhxOuBeDykZy
OHhdd49EYxWciTopSIM97XO+Vj2Z6gXZvhnTVC/S8b6DFNuYvrPtdbO556rxG49z
8ByaHx3pvPygSsi4eyZy4Ff9ABCL7tJpjiMYTiNF89PL3pGz0Q9YUtocYbut4c0c
0bFVjaauj/Lt2Jy/LOGAS9F5tZ1U9IRzKjleW25/KEDjijw+p+Gnp47vwg0QsrPc
ReFgkyfOvvAFxiAcKEXalMj9CxEuLPSazM5frhtvTMbaVP8TcubGQ3oD8HG3J0PI
uClufwkJPUDhKxzIxgCWvOBlIUXKJ1mTla+WoSJ4RcW7G3Rr5wI/P+ymwq33Md5A
JQtX9rB5dbzgqIniI77UPiBlqi+GwytAqHZCh+r5A4UNdCISqVjtp6lYWVAqiu4X
+dHuolq35RlDixmL2CfEL6b6iwfPC5BYr+56wh4wE7GBxNmM8IrOyZulPKRDQH2e
mVRikgYrDD46fveMVPNOVczFByJp2237X8ITOVVJJNnBDJf/uFr78Sj7K5IS+hOb
D/A1gjiC21R2FFy4joVZBL7tYMG959QVGD7f3AyEPVE2xCpUz1p92PvpteaaNCso
pLaDwMdZx7w/IAsLhWv2Fz5/N7xU02CqjzIW+vlDkzmBYWRc5a9+GRMwG+XYBRcl
UxiX6Hgsm48mKugNDi34c8c0Bc1W/4MqrL4QBNMps5yYH+gbvUnK2ZpqZtIF0kwY
ysgNjq8+Suke03QfjM0yOHZboQ9jkYhHbKajCNDUMtZMFvEjnbz26D/Tt93+2uWv
hmFPo3+Lda8P0zIVWZMhdL+auGKvUq4+ob7wNJDEivjBniuQQz4dh70zro/iPy+/
8cOkR126BukBrbB2gKvcJngxwsX6JHYFhDvmQ+yiTlx5ykarnTRf5CV3D0rNDpzi
EhtPeyNnI30AfNbzG5Y05l6qMT8tkleFqdhCSVDTCpMdsKvuvVU3xtda8VDCMS8r
5og9R0NdURumpFU4z3xH17DRY6s4FQgabsQNvs8ANNdoySKabZD44OwDY5ZVXSQJ
5wNiYi1otH2QWtniahCw/BvE8tUiLCqMXPtvqGlKhHpcK2fBtmby7Hl5Y5bCUH0o
fKTfkzfFNjN7vuR9VVKvQ/iydCfy/L6Eum7fRf1KoDDoCWb2ifCNlXxFHSWpGd5N
EM6dmpEUUDM6w3csrRHuv+mcC9mrkzUp9/KXNUQxBa/JxAio4jeDG8XU/lZiYJVS
N9bSz7WK60+N6HGYAUOWCmmGGwx2nlM5FYagY1+D9broK9hZ7tY5FCFp1mUEon7j
P5elegLBn7qr9QsA3m2GQQADnX4W7kKw5gXH7czCqrSIsDNPjojHMEn0M64GXuDq
V9Rj9bsGPzJtF8qc5I+ZkZPu7wQniwSSSIHFMo+4IxXPfqBpoKPfYk+vqlng0FEZ
FpwRuuw3NuG7U9mp8w+sMUzJmE6C/1W0qA/xX2lEpMtaEw5sMc4I+9qc6uy3qCTT
5zSGScrKR+Vll+0Cum5+73ZHjynMcRciy4+o+lnST+HSLlBodq33yFsk5c8MdAg4
012ZlS/BHZyp3z9bpJPgWCcOTJ3kpOWgwbq982bDEWsKmHXnRdJcF1jJMWanjiDB
GyQR6TyiaoGQHQ6U3VC6gF1CJGBV0pB0qjSxZvo5WutIkAwZDL0guk9dGga5FYIU
8mFRuKZqTVslNI/NWmrNkdRQfI1wmtgHZHyRUxtlaHj6eAhjPzhNBWzFwVcOS9A0
y2uuhyU3LVPHwi7acOf6dP7vUaff/sPox3qFbzHMIpaAQz4lymy9voCWKtwjxfbh
/9dv5g37Q36m5smAzxr0MV0odWLtFfkiqR8UIyTsYUMxppuYylfoEaA95NfrC/hp
7dqhpfluZ0bRNrcAGALLMHAFOEq08bUJ7piul3QH0VoBqo0pBe6GwiPkfkvRjoGN
9MZ2A0rho82lZgu2zXYRhfRT5jDbgcWIWpXNUOmZte1Vp4Q/dxQ7Qw9QnF683Uox
rVSCck4DYv3F8T8G6MPT3xmcOZJ8tUAZMIW5sge04mi7fKMoOOqKCgRutZPFJvgy
UQBR9/kEzgYHmeO1aXmo997RTySPDQRIXg/5VzQSNpMdDRnlQ5xKcoaU1xQnwMEK
5BJImF6HR/5Z64ssSTEUqhGqFtWbAUXnbSZlrd0uJ+XsMYUM/lbDwynklX0VwHEO
DmYQjqHFV0LTVNd9vTZO0lh5v1i7yZR+INDqEb4diifaBuk15duueB2xC0IbaJbC
ZmIdwXYPCKwmFOXz8IjWU/p/1/9MmLvIevqc1cOwR2mApfBXuH8vwDMuG2IkkI8a
HRBGqjNfNFvKuKK01/SvoJKUO9GAHu41Qtj5ROq5uEMi6ZTx1+3/S3cqln886+sP
95h8BF3KqEwf4KseRX9/RmTgHlzj/Q12mVZIRjugSte093OYgzN0yo0K6xwMVfS1
UzmZ3+jx62YWwgfuP4QO7alPysr6rON3jWHJQJWY5nu/5UMTw8Wb3MVwGcLAkQh/
tg7KcSy4ki0NnPFgnPoD7Qxnp37bImmkOH65UF1aOq27tpw99p6Q7M5IPcxaxdrn
BRMnwyT1zPVVhP7yTJqrYoZHcChNYODc+bcQK3O+RIuRN7wkro5I0E9LCHBAV4BU
s5vdzTadZue814ssR7LzkDyMK9lxVieOU31/BSP+Q4inZEnTcZx5ipz+4djybp6G
TnggDqBeUubuk55VQ/FjPgijn2do3xAgLeYhoJYUneagczogogMSNVuhEv8mJtLX
JkbVfCbUr7HbAZlprhm8ubE2lCm9Dl8Iyx/GE7ckujgwsdWPLCMz3cOfahq+mC+9
7xyqe2O15kOgS2N+PEDcGzOIXxBueWHzblaoo5osXTyoLSl8kA+TfXgb/5GBQvHx
gb5i7E1AQmkPkT1AfT3pUNKwBIu5zpZJqRJz9TqEymqnwjorr6TrCxtGC5YXoRaE
4OuuWtdzP5+JXH//hJaRKpCwjHNX14Nqatek22k8fNXhEGx+YbgFIl+L/Icm61EJ
zxTRCmThOYP6S6LfUp6NAveeygsgHJnjwWrDdF/lkGwXya49YTwk5oWhKg6QJTJx
RaJLJ5Hxy/FmZcJ96ONaJe23i2U3ir3BzoYkFY68wtLK0k1CE11H18jxOOsiNQA2
T2+gZA3ZyIDCOaVsSomEBGZEYzkeznuqkxWq/T44UdNfhOuruIHas0XkTdcKGfDq
Dl8DYo+c6CcMAUUBUaJwdN/2m9Lzuf5JW2IQzcYfhv5sKjnT0UCWw9T2fpOeY3KD
uGkZ0kvat3iJHAYjguA04gQ/skiy2EWrJqZz5j/t34IbdPPWVk45U55ChwxwwjOx
yZMkBL4xoits+D4Zcr5PNzC99Iw86WzWl0ozySRCef6fA2yRrfcni5KWvzj4djLv
YGbnGa/Bqvkx/fAY8t0gWKmw9+U7ZFu/XwH8sNu+V9L/wJv6+l9W2j/Bt/aHWaIV
tCdMSLn5teuLOXC8Mer8t4/eoVqJXy4GfvlwBmfzB0WMKaJpoygWU5DNBMShZuSg
nBoGnTm2mhD0VmQVwCO6jaIIrD5GpnMhlcy1LBKn03QTp+p2llOLMeF7GZoRWIJU
VVbkkTCDjyW7F8W+jP8/3hXo8YlCXgaUr8gsdCEHLF0FxBuDHSFG00lpz9gSRp/i
ePBU9Pe7GsMW9uSIZ1t1UykPawdBhS25ptcTVO2r+lh69vUZmfNeGYOoKJ9bR3mf
sLQNjP4+Rkr5oStiadGbthgFJDrwzVEE3lHblYDe7I3s7sDMn5x9+41t2J9TUsWL
A8iPjH7hnUQCypBCGsv91qv7s2/QG9EV4q3yoQ6h/eN6Xij340xCVUAv1MD/K0fe
C6AhHVexHdmKnnvkK/Pc7J6z1YuFUNUsVZOQmkXC1uM0grfFDiQ8face9qMGYoSB
RdS1W2Ja2BF4hlMFykP5x1P5AzwVBmmGTlPHRPfM6WfICwpB/g6UTlnQX7u2bT8G
FAiNnsY0pnxztZvdwGEmOqFL5j8BANhYSj0CUcYXR9Sacdvlrim5CYxHGT2c9+jJ
z/U1V+eordkPitFCS5IHMtMIX3eEoX8JzHq6zUyCk2Kv38Ghe31R4UCMgLEfFyRX
9mZFYL3n2NbrdMsuhDtEmSy7ZOhyE95qd9/qhPxrvM34xLh5ZT5DIf72KrVwVwgc
hntTs8Mq8blC9RsiYKY6pTdLgeyM4LDbvq93MAafJ2OpjXTJD7D5lryf7lsUkcrY
VSvJFUQDqqLQW4Lnkldyr74ttozHKndKy+dpKzKGKS5oWLh0Ao7+FoOUVSiVqPVY
3LDb/NwcGhwYtakumAOvjwFHGd9T+Ynz2YGieaVHWs/Nu2eZ3ZrDhnG/i3+41Ur5
pTeEeNaBbNFFQWDF28FbF7IukzxBA5tZnMcOrmTJ3UUZFey1oibNGlcAFgPK4QlS
GTx0756gfTfTSNdN6ybGqGTMfYglohw2wyQbZLXyYuSvLmfxStmJXas5IQtgK5sx
9NkipKjDtyl4mjKhc8fNIZehA3AjmbRkD76ByhhsxFrM/PN+/kg5gxezV1IoviI6
7QcK1rjNCM2sVOX0+LJ+rcrKwmqZfvGgGRd4gaKZ/8IhWIgWgA5jWB0Bi39ZnkSA
08YxiiegNECeWVyftbFFGtV1XJi+OneV5HkSKdDgysZwz8Te1kEF4i5pQv9OBvj5
zBIh6R5tBQhI1148FHUy3I4e6JdVS1R7vYmvllAuo4heXciODOPElMBVAvXvuKg1
AUQBFaJm7I8Rb1KpKGPVN2SkHsE6YC1SyH61CdrBkpj5mSe/XpkmiPM4rbCya2dK
tQRbLKip6k5GW9dPrWCommuvRSvIoAmwKJaTeh7V0I/p/j2em0KI12r/WIGQajOH
047hnxwBE20WTOLqSUgvfuzv8sIHKzQHZAd9J1lWjuxK6sE5dBHEJGfNYBTfgM3s
rrAfDgsW3a1RGAQjnTJHTl6kc/kFOdsHaellvyl85Qj8yITlr6/YIiwRsXXz/BLq
LT/nlwM6X6OT0Uam/QNncCePH1wnxDp6l2h/DzQylKNReGLrIwNCy5Gvs7wFfGoE
9sJsQ1iNXnI9Rat5jMKBHzj7E9aEiphnuZsJibJxk0lDHLyxzElf1zt0I38luJkP
eUSDbXO5C1g+nX7wCJZY0wWFlaE7W+yKSiApMCaDuWJjveJYXJiem/CeDHxwiBJo
pttoSwkDjueEYJmJCWcgZqhTN06XGAeew6P4t+TC1vQ2XzU+4uUnAzQ+WGEKqtde
MoTeHnwHDl+LOCtL+n/SVsQGGj6brcxIPWM4e6qX4iWn2gr+qcWusnYWEGTj6I6g
KY3DRCtQg2uJYYZ2YK7G4UJyTd2PCc/2QXl6U/CZGHwDfK86eNn925kfz1W5Bmpf
s+qQb2mJ8uJ15SYF682sAqZBlx90HXlV5vernHk3kxnVKTfawdAHKGtXJrPqHooe
2/GSCAM7z8KSoT0NJzJ0oezjr3TNyXQb+yTUClIxJp4nkOC+AZ1piw/PfbuZHyR2
UhfwhU+PSY+kQkBeDGKzuTA515R4wTqjg5nqWdS69vT2KB0oQ6UbRhucm1lX1Wnl
8Lk9zn55eJowEo/0QMFn+aNFzLeDOin7F8+9D1BlbreL4S5texBl0o3Sp0BxJhCq
jXTcHNuT/Xc9VPmsCLXz89LPpqGt0dM/ynRzYl+BalIzNICzpUMtcfe6kAr8AQAq
R8WzYKKDys+3tW2JdBTUKhXzM2qnY22rwkvf3Nu5e2dgQHdvZmBOjobo717DtrI8
EaSjE+Vzm0QtR+csO+DmVUjcwXA/a7+mxopaVK3BFqa8vlGNAfqgB+sIQOrUSz6m
pkznXgkWjE07YzvxFrcQdfDSn6CRWN7BiUb3bu+AmWc3NOs7O2abXprGlQqY/RDQ
GC5ourQfCAHPPzEQzTp7gfbR7AfSWapM/ZyliOB+KrjGh3gnEK9q8D9hHCtDDo5h
kJhisYYpvU2EzjEPbK+mM/+lFI00A9f6rwWi4ca3Adun8z29Qz3G7k7on3RcQbxV
wG8iPsZ6kj4qmhHLmlOGV/zcK2w3CxbjAWf2mXq5usPLZjlcJMZpBdLNRoMeIZfL
4jk4fGOo5pXUaM2vkqwUZmktX7zw+87UdMmC8DsiwAz7G+4g6okz2zPd/mjcJJzP
/YPVY8qlwjiVN5nswZH9DqSdNPdv3cp0jBRvh6IpapUy42OE9lMmBxDtISfHUHJW
Kn3mUYacSB+of0fbAlRSquCMpbt6kKtKvQmoutOFUtxY/rnq3vGgQ7xBlx4KzOus
nlT1BsonDw8AJ1ue09FtxSFl6FIqd3gXCLbHCKNOO8VNOIqwSqhvPt4k58vAruWv
tm7B8luZ+QKt9yXt39MtHr5GyJsdsmb42T8WKtPiekA5asF4m1nmJEfQw5h2smrY
uJvCFS3ESsaOnl4Pc3mfISjP5DAOniiKzZFl0Jb920djujVYCjxbd30VLBGCQd2o
JzkJjlDD6zhmGTpXgKlGBZAwMdfjKqLqMHv4ZgOALiia1nkPonpg18iCeGUI9sYJ
Gr1nTa/rhhxtCntM13gISSncGwWiTtrVzy42p0AkKl+p0DA0GqZIi74uBylF53iw
mzQ3W6Rt9CXVtHfi57cK4nYMlhl7l321UDo51dK/M8/3WwATnsMnunKwQIBjA2eX
CzcPJolqNgRlXwW8NXf0e55rn3ScnfCarrX313NYEubPE3du7ncgf3l7nImDSYAa
xpClk2YEuED9y1cwT6Ng1X45mZjimZbQWcwoUOJS53PYplLGvoufBnhM2tzKcmmi
s4XpDZ5CzNALJguPJLleLrQiZrkfcsAZcGY3ejaSFEAs9qzwPzWYPMep3+r6tPk0
YwsWSOEMmYZx+Ypyx8ZxSihhWfqn+dVRY24fn9nFx882qhm06tfb5O6kSlv6rlBK
z6e9jbtIIck1r73Ds5ipwEIMN/AuqxCJJALeH3AhB90FeEcutg7/1eA3njcESAS9
U0Zqhe20LMd6ugggtMV1Y6thktLWrw3Nsemn2JAiMwt5jybZSZ4VfwLqijB643E+
EML4U8GhunT4IEsHl2eGpl6uAEWI+ePugfmY5X/jORWQq1Yr0NN7CPEPHFf9H/G2
U1jyKNWs7mPK+t1GbxljO+Vx9/LBiVHXpPTV2dNmXItwvbR7W/KKLTBaic9vhCwy
Pus/sJDrKiSSfVH5UjKX1Op9C13JNdoBWfP8jknF99vch/306qPXjvTsURN62NCu
qr694O0YPNK0c1iOUP0OZagrLUXlPmtLDkYGxFwoAa3b+KMEGf0SFrC7YQe5B8NA
ZEn4Sw4UmabntSuM9bLw6d7XDnNZ7dWnRZizvdqO51QZnL5V/+CN7wuJ9q01BaFl
C0Jhl20m65RsGLQ2dVSmhfGvTQQbm3172AiSD8WroHJZARNlT3F3X83GXriKwZ2w
wuXldP0K7SMiT6MnVlA9a8J39W+PTE4HBmIM8k3CSbHKo3zFxJ7CAVVOuqGcdM2t
5tw+X7yUuUNI8wBqKuTgaj373mXhRFDlzQ9P5ExEqhtbfui+IYOXWJ6LHqTX90a1
dBZYEd6WtK3QWrzGDXeJDp2mpjduV7XuHMxLAkTAIwVnnNGBvHdHO9o9lzUL7nlJ
4hXrI9m/EOvyI56iM+7UeX0UW7l9IbnodGE9LBfzWGD0Da4AZFfanHrMlEol33pN
cMYvtgW8C9hx/qvx1P5VRyXEuYIJqq/UUsZVH6bh2vJhMoKBWcqHdWMIDX3dahPg
Kn2t54hdHE2OJz4E0yYDJpFQ51YUvDvfgELasBS7dWSa97g+8fykJsNQj1kEfi0S
Mjvs+bzbqA2xja+YpsCPd06tsyHn2OG/+ABe0H4NJh0upTMEy7dGbb4A4oMuCXz7
0qGCknp60ualJKMGfa9EMJEwyxFkyS99cv7mSxWKBq6plOU6WYnb6TNgVhbhXaOJ
XFhjpopq61vMGM6IB9RVBgXciyrnitnhY7JeowljIA1B1D5xO176CoQ3Il8SbQBB
/gXVdq/0PZZ/gyBw54yE0A3OQJEaOsD/+oJVOd3JsUR9V5jdoIj4xZPvL+RGjzrW
gEwIaZDyBwarHb+/B7EMatsSVHz4XgPgOzg2kGKg7AAUzY25CV4ZIcoOVTyRMGF0
VmO21OGUBxJCBjhV0cpHU/WbhiZS661rSKKysEfWkFwbnHd8nlwi9/Op2j5+t/r1
ihomEJBCyfkuQ/m5o/t1e0vKV+Ey3ynNogvW3+WfLxkPwR2Gp4v4VICjA2JW/zZ7
jq6qHfa8rOgEvm3OL2afRoENTVuMt64ySgv+yYj2UiA1u6558qFud+VpAnQGx5A7
E3tvHBH1yDihCWu9qdlJ1nUZmVBgA2B7WPF4dQ9gVjQd6JzSn1RIPLQzkjefLXLM
bG5NR6s6QweGzysSX1qX5XJLoPXWTdgkfSSu+34wndRrXqiXozlQkzojtbxsBfl0
ZYIH7g68glm59M1TdZyvts3mP00bAc5BncAMEMO6CzifdZN/KXpHssJYE7k8rJOA
eIC7+9fTNNjLZNp1M0jhXQcCVZ2ujZYpyWdz2OL1TMQcr5QNhFll3pSmBr24P15p
D2virv4kJIR+sYtXLWWJlkoQBETJXSksV0vrmqGDaTCS6QGu7BaOH14I0HAJi85Q
i56BLyD2QQZU/tUfzbOggK6KpPcKO6qYgRSkYBJt1sra7HJH/OAVM+pi9Jy0e4nR
5A58/tERl6qB0ck5FUoFDKTLXgFJzaTqfZ9D+SuADEBaOeGyfaOg7Wzx9BA6/sIp
kzxArnlTyH+V7YrJftXMwqCkZmOflD64N7hjc1+o3NFBumiILNWAq7sey3cwgoUw
LcpQQr7s8hALWgnQvHi6h0Z8kVK97DslMvPPza13jsrhOYAhKDuCbC5ZOJWqDwGh
xn+1U29x68tvkrkuRLVnDhwFBouNmwKZVFbXCYfBk4LRmxow2J+eB0MhPu9JwL4F
6YGYYyXnptTXKbpcYIMjlI5IkGnBo1FSezttN0aht6JINXghp5kFD9yLrV8/hMvn
tnt5hkzfuR/A1Fk/mHAaPWvHyDT1I8k/Rs7ZmLF+NcXcz2kXickuOMDMAD/nXvHW
U5L5GEYUPzqQHLBtFDwO7XWQ0jnpWAijXSeXE+doiv9bICFBel4p3DJ9IuSBXF4D
nhOxBWuAcqP/c94y1J7YgKbcHHk5sfZ04a5+/KCFMFJCeqnFxiNr1r7GdHWgCrNr
xkP9wDdwJ5yLq5tyQBtSSxArLoJQKvIIqJcxSGeoltPgjFzaXCzs2uUTEiO6L8KJ
Gb3OtGEgdDAT7EpnpwiEe9h8Kpys0e5SW9ifjqe5jfhXg463SrmOyd0FEuuHcXLC
l1wUB9x5ESZz8m4EKWihkXjaa96YSSoVgYwEH7eRhRnC/i8+KV9wUfgY8JMzB1Gj
gLn5Ww/vNMu2smRu/5Z9aGMgkUpL2SnkCjhvk7s3XAMi3EJT9ThwLfRfyMvQHRk4
O9egvegfaypie8FryLq8Ea/WZ9/sjN+BKe6hQKD6khoKIdKLrcDYgTOE7T2qCDrb
il8pN/nw3eOvP8sTohCV/D3GnWlw3mC6/MMmatQi9LAGuVewQCyqhf9v4fqBST9h
cMN4uf5AtloDOkJnTWB+POwIIM1+9DjEW7ykjXRrjqFDbGA6TYXo3L8zckYZDlHS
o3XWUog6dcOmfDKz8BuKdUZcWdXVf4svJrSxCLDRzAH5vf0V+2KnNByx9mGSUhKa
Yz360oXou3oJkVDHbuR9D989fD7SzEo/l5UVaMxTvAsZdJWRc0LmxECOQDEbUJUr
VNQWd7FfFdHp3BNRpNpbDCRSTRWYZdKKeIAJNrGooP+TdSqAZ7TvWdGpD8zYodj1
ormwpHlYS2uh1bEbvD1YVI7vQoozsY6N7VrGXRFFUXbIVsAVynFjdddi0CzZfua5
ua+iIKEQAMTvVTyM92eyIeW6dSy/jInuAG6kq6UlDr+tB3AFY5qRtck5k9G11fkR
8H1COvH53baLL4FAd0n6qZhd/0Dce74ZYWLzFaRJ49GxpF5gdxzxEFgWzlBVwmrF
BR2kmzHCCiqrmUOdIG/af1pL1ZpF0mVHri+Zk3mkq4IpSRU0z2+aS4vhg9AwsF76
cC9Yq9NsVgMbVqY8gqyngLAaJch071Z1zwtvbFiMuJwgEjeya7p7JCKxanlG8TBU
JdBaRZqNn3d5D60yzePGWZLOoIy/tNboqXsH3T78Znc0uyTXZ3Eu1WpV06gtQkua
3TSejMic2ldVsZlLfgVoPXYOSns2zTNY7J/lezNRtTc0NJ0BQf7itz1uGEC9+W0N
jfPa6ehklBq5KQeWKTc36fG8s/ETsSwm7+yZMbkIytfiARQiYMY4r6oky55NSZ7q
8EFSWPmdaGuFqKpiUgPdzEMcsWHLMUY3SqtDHSoW+2Nyvv753GUR2N6xjzdjB4Qa
R+YfA9LbkJWx+mL6Y2Xiti38NPHcetWdYV7WPVAF3BKxQHQE+u+/Rafc0QbqyGKJ
ZauuLbGw79bsn2IIdIuWUVASyrcQDrIrk6aPv4x6wgJkKBEcw3xwR0btnVCsPtqe
XwL5/MQR8KN+wj6rFtfKvmGsVvMjtyDrvOMZn1p5wClxQQ8ZhHAeHcG2ZDMSABSD
tyiGcFDA/hq+kXlc/qqTBYevPsgehM7e8+szw3BOLvRqQ5DdIHxUGFTtHKk1r5PI
Q2wCi4BrUpFTk/J3UpL7I8i+vsCMKcSVdd3sgwcJADkFF635XSfvrkQwYN3mAPEJ
2PrPHVKgZBbrbHSmJRQy+XMh7lxJM/ldFVyUBD563C+WRQ/n0L2j/h44LAaitMwC
oFcjemNZszGgxwXBx8niMa8E9F31UbhkHTif9kVVSBHFx6OVy4hrLFLJVowHlO4e
8YE4u9nzM7TahvAgwr1YjlKqLAwh33IQrEm8nmW3gbyjAmOvNZsmD/hgXibN/A/q
8rsKFD3PIQMgy+T2B11Ra9YmneTJ+YKtaywteYA733U07F7cbraPrB9WLPyPADc8
OY1q9vOw7I+wdggy2POZc+tY1+cs/3VvvEEPnZTTNS3pkOnNqkf0pF+h+ep7Hk6E
YPDci0KAF8TdN6/fm9BKWOPg+ZWKHaZqoBR6FytujGlSLaZN7oPTdgZrS37BwfKv
840O0XY/Cddj5ftjk1u8d0v0qfU0EPYLxVVu6hbI0buVegtY27WIwxzFo/pftTfW
y2WJ6bDukNnn/OzksAxui94DBZOZfIhB7RO7q2fz1K43Wzx/kLC6tc54f6GY9LPX
IFnU29B98JWyqoLkyPwEzAoPs0THxJPf6Y5FMC5l9k3bPKR0fCTjkyFqfzmMNwt3
tGkiWJVc/0Y66zgKejHnOgRR7/uCFkGDPZiVEEl+jVM53NiopmMjurb2tUYkLMtA
RpZ7pVRA6xAP/liZ7b0kOWOjOKHGVJMl/XG2oSWpPh3xCqXCVmV8xFRofDLcjQZE
ZAzsM2EUgrTIaj8aN+ZKThkaxHHupNHRZOU+3oCzS4PQKgK9eXRibFZYPT25wbXt
LTf4c+z6gBIx8eQdYINp4nZAo2wakYQymarHrmnun6fe0lVotoQce8u1LMAell3b
TXDK0a3+XEOwtRmt9v6lm7N9M/M7tuCVgzLY+bG2KKqx0mUt9lyd0yMM4SpeWR6f
QY5v1ITxJZ/cdJ7uN5CzJ0TkgI3WmVIGE5yw3BED/cWrAi7WEgOOzmu7oWrpeOX7
AY7kUqXI5WhQBw7I4AYtazNWvnUz2oUzGRgFhLQb+bLk6DlxSamp0evEoItXMC72
sjB9fQPH47xrUi+Oyff6XmL0SLVgLPK+BZySZD2Q0z4a/R/Jm56jYhIiPEgk7aAG
uBF1kWbFiotQNqNos3jnt67Optk5lC20w+kPaGX3GTdwroP8RqJSC06NvXyVPu8y
rkFVVtcY12RdoNM/uLM6OymwN295CFADD9+olpQprzjS3i0kxDcVMonWPCdKk5KR
O9ZJnFrfgSSA7ams6W20WxcvrSJizRl19Uj+PGPJ8MqXumscWqtxTkMSfTAbOOBc
6lXn9NyZYmPcabH+2rA+qnBCEuBADmOsu7UNqm1rnHHTzRMdStnrjoXPvbFfP1pa
u25lXoRD3DRmdF7+8QfADiM3PfGOyuVurnH+9GRr04gcAP1XbSBGcPOEeHsgk84a
4VIywRK5vSofGu24TQrp8Pz43ePlm5DOp0ok77Yvc9XoHr42L372GHGFRi4QqhGa
5SFZ/TeBeMRSEy9ga4wt3fygh02MXajobdrcXNnVSHhA1XI9y8UViXHAlPvhaC+e
LWCmC+iECmvckHT5O6AfqGCq9yy9vkD9SRWlteZlRzG/fN8d8pi0VsB3xybv/4Pj
ux97aZ0U6HEm8MQllCCTI4xCPaBA08dmpWG5QotBY9SSoCSnDWWNVbJM14TPvZ29
akNRaoTwbVOJk6vrPCuZrgfZDP4GICMxkyFRNXWpHghrmf0Jv8Z//sjWR0fKExAd
teV2iSdKHtbzWYyoQmNgBLLS0bUm84IlV2dKlkP8BTbvGguh2dVIZPc5JbMPsd3K
kIsNFPQs5ne8IG4DvMI04Y6a/T/6YmTVGfxZyyiK27Jmwn+in67CENdXjGpYYBup
8Y7/0idu7vrcg9rj3uIjuGZoDImr79wzZPTSXAQz+0Fn545+eWawfV/gc3pDdblC
VYE/tB+4S32X2KybOPuF7uBFYDnkZT1osgdfPmVD24oe+HAzAhj18asHA0r1aAvo
GtUrpTwE5V0UQI3sJSeZuwk7MaHpYlX33/PUMpErqfYgSvnBON6VEcfomiAhfZ97
veqmM4dEDg090BdUbpbKB4kV84OY29Gc9kJT2xtZNLTRNzlloFO64DNiTzhr5HMw
tUGFZ1zcn5ZTD7iPesnwQgvg9dUaeamJMqYR5VN2ilyYA7VFl6H3o+SwgU94Sh3W
UbTUiu07vBQtG0rXGpP+xdJ5GAoQ/BhQS3xavKiLfZLLCe7aDVuQh19gP758YPDV
lQn/G4CLhmhWAEa4ghOX77ERWqGx25SRoMa49IIaUXIkP7iyU2JBySLdZE4QRBI7
sGHaHFLr+DveSwU6FI5+6FNbcst8nyMH/Hqw7bQf3QpJN5WqrJ3bqHa6ohgdcC9B
Cfv41rUj51/pKUmeK3gpasIuXgHbitNXQA4ZoRQZD3WSq8ginUPX1MBtRmKbRy/i
T1+vUaHdQYVLYmpt1HbjXhl0PUXoyFIaj6Jt994f0FslOOKEGPMjgaa0E+2qXiXG
78XLR9moutF1EM05lsgYI96MCZkS7dUvJX18/GV9K0O1cxLh8gU7V4Ds5+HtbwlY
js9n9IWnXDgbX8QYRQ5oe28HN8v0OUb8ubemKs3DGKcpk00Pgr/xPiWxbxyYaG/X
SC2UEBrz65rl9Ww0QatsOsO7MOLJviK2bIliWXygttkfaedI2JxfhVECI3sOj3sv
BjNcthAbqTnKZUf1JnAXc85M5bt+L3sYJtdfi7tj2NyDCtr2w6hyAyoFdGkBeolL
DVkx5BSlZWtgqkLEBiyY1yPzwNXVa5sjx79PICNjiCfk9nxRBxBmZyOjicMo12yS
QAX0dWNlXjlw6EOuLzShLvxQMZlNpDeoD47b+6Ka3ni2IDAO3XIiKAazc/81JenD
6veaNpdIUbJzwvNL+o3xI/xlKXSSRKcIr9XwJS+lmQXNZb/mE+V83E3h3g+dCC4c
P9kKEDKB9dUrk7reYdrGQQfVp5fmceECBaxUcyDyLNCR7mXSAqrmZubhyD0BWxua
t3iE1svTjkFmXRR2sIrWpsCh4+5qIin/Hir6eIrQprEGlBA5AGUysJruEV/Ot+F8
PAvE9Ihdy7b/AKUry6tDUtKeUX5uOQogFw5PTnDLkuUweUYbEiJUUyNw1VtKUsg2
ot3FSnHAhE9ggluHE9rAVUaDsv1Rt5LfK/w+733ZHxX0aSbdJpgPgAR2aQuoUaxR
ZTNkW6a6XNP+ITT6HhzPTaYzOMKh5NkS+gAWF1uGZ6cTh21yO4Zc6vHV1Ml5RoTU
PoTMGOHt/TwArScmArb0Uq64zxRVRyCM998xGqJ0cLS15mrOL6zoUmulsBQyvkXy
smmNu0uzvLS6L0nY8lQ1gX69mpFPBmf2BONMYLAP+T2ZDuuGIn2TkVmGqdvnZvvM
mh2gTPPvAyHlFrcuMyTk7jwws21jXJbEkqUTbYIgrbE7H/X7X8DuiyZQC9+//072
gwwIoD9xBn8xWPhoL/KuTNLZIJMzThNBB8d8qt/1fwyEDQ4k/MLKqxQiZBT2RC7o
DCRBEkTHbCZuAcfQl4+U68FOwC57AdpU91Wf3EwMwhFxY2RRNjbrZoAdsIpXNmUm
MAr2newmjhNWi6WKJVbEtwtZUqKtyWs7YrKvNrdlfBzsv5fzfa3y6Xwn4X5vbUm/
xOjlqGf0BXZVW3aWJgzQTJYR4/aLlO5uL+UTlE+vxj9/wQBrhiPJHf93FqLMPyyE
1WJ6EZPxIoI9zzYEQPTwYyS9J3OOZ67QXzJoStwssel7JF+rLHXIyGPorvhNR1qt
96kOhSpGg0ZgMbqY6jCxbLexO1kM731IbLsoaOAffdFLcCfc87tMlXq0thF4dGMw
6NOELc5upIq5rykz0IsaxPx+dBCoYKwlcpF0K1CeUv0yV+GVtF3GCBLAWO5M4Yop
wz4R4ZqkU6izg2tREnmZHdBHu/m5nlESK/SQmwO/JjgiB0enXnlCBs/L3af0hutc
Afg6UwEo+ACLl+g+YnA19UUkwHFa2Y9WGAcw0piIUzMLSu710jxI7fqWa8EVZ55Q
7c46IcwzpNIBirfouG2sQAmarKCx7aXFptE3J3FRqL1t04qI9Tn+UHZaiB9434F1
txUQdU0V6QqETVgyjY7EM4Zf3atiSQvhXhT/siHAaWz1qtMeVjZWMvvfv0ISEy6S
IuFk9ALpKATS8X+uG5F277tiWfbSsqDi9m/bI+KdPjNK0C6UbR8kBPlMW6atQ/ob
F9MwGLa5sp2V5wKnwQrlzpr0uhwK9KLXcxEjCqD2caNa6L3B4ffceiyFI9lMWJZK
5UJA8LZyeQZQorqoJU4vyXmp6lYfVlEn7UEQJwIjyYlvojateBGSCAAOlRrThcV+
zlLlUaDXdc28eUAcW0pVrtwJoiW4xnIQSm0gR64Evba6nYVmNkWdCUWrty7+AGLj
ILK71HmnOjDhDQqTZXG0wq1mPXUBCkttyv+2lVJO+aAUwX8beQKM/mbvgQyOBNzY
RvEHbMkW5E1+oSJRfOVCn3WNEPzUWeOKcqXuemJYg764XFclWDX/5VGo3+ctUXVz
uGPsz8AH5N/Gc2bSDECJ3s2XQUbnkK8qzvPrSqM0uNd6FvxVSfBTYkGVhqU1V6lH
dQ7FoXQG2PqXPJItWoFuhzqiipyyZDoCBpU5ROIKNWserk+Lm9hpUdT+KmTnFLqa
ZNZscMGi0eBrKQSpc5DIPfxLrxs1CXlylxCk5gO9Nor9Z82FMCcv79aqs7UAfebO
fM/taQH6+TmAGXm83x1l2URI/Dm39m65/Mp3+/iolnF8URCZqGayQZTRqBYGUmr3
JkNOXJ4y//LN9l+Pz6MN6s1QbYv6xvp8x8jrOauCRF0RPrlWjTMcspwBVJ7A06CO
fBYc5HG/ouTpB3REtg3N3e2qYAjyCrDjpJ1p74X706SoUefj/FLDhKNJWw8SnUVz
Tmzpxe+yqOAjY0DALRYhV0TKmtY5scp6Lnn7TAtqngKzD3Y/iArwtq4gX2SqE9VR
2vfv3JOuJ4C9hvYBzObz4aiKZeX63JFMigP1MPP+tb7H6CIfRXDYsaLa+m7bg3Hz
CwbdT8Cs9yKdflVdvA5CK+4+6MDJOjp+YJZoi8RedDI0UWYP0S7omjddCYw1ozkf
MsTariTXbLJDX21b0C7IKZuca+Oz19yQqaVzmPHt3+EdxYRBSa3+aFWl+UiaaDyN
khsiBFg9flSC7WjUfcEnl4/R3eVJ03ov5c47vuKaplDrdhpcYCFADO0iOP8HvH9I
4HOQbgWGHtLPK08n7F/oCKpWc9maW91qBC3zTXdv6BbEifVe3zj3g9738wakJlrb
rTJzMbF0LZB0yX6Hhv1GedT5mQfEMtsHO0UO+W7SElYYYpiU9f5IyJWVt3fllZLX
usu0FNSWtHey7vivBLD/MvwOgcIkJOapZQyVBC9VcfD3zjXvuf293kDJmG+Rf8pj
T2i2PojDgTUt2YQUf5wqLqk8iXJJQMJlIfyhcgYI0PVwUIRlxRiCF17DjTfuA3JK
t7Ql/+O76a9MsIRRrJuzjGsMpc2bTAoNKc7DWrZ1Bo9hll6WeLM4SnfXlu19QHw6
D8G1Zt3BNNIpspzu3KzMaz88HUc2dfN58nskg12An6SOrzKLOtBJ+V5s19hlyVDv
4/jln5kagIJDVLtSAj1C6Rm1i6uOqIf2oGTPo497zmZC5XPo94fWUUtSmThqsv9n
PrVQQRN2oZjCIacUeFY5aUKrK1pqun0C5ZDs4mik27KVW7STTz4h97QJkw4Y8vvu
0USytYY/HKXzF3+u9oo2gQYGiBT/FdMxlDjXGK1F7bF7bVDfNW8Ui+jx4or5lEwe
1iMQUhe85g8tMZCO0KZV9zcKLp/RihchPUoezNHyutO/I7xPl+X7I8l9MEdTsruE
2PCi7Xr0ZdD55CkKv/VP0h4CAQChNxIfjOc0FoC0051hvILpAdr4jC3lu4YgWI7D
OGSyhiL2+ZhYr8agat5e2WRPiwAHS0F6xVH+/Q75c1W3JvG/+QPZI2eR7iz0X45s
slxbjZL24BC5jJctM3yh3b7w4e//pvMC6pUOjPePLSSHpIZTp6S9W2NJ5hOuEdhZ
QMigA94Fv7vivhQXmU2gA4huX62uj7Zbn+uvZfHQKU1781Dome+cwVRzZegrRa1f
ragOlD667pcCjTClcULV5z6e0kTgvO9bGXz+o0ie3GiR2fOerrICJFiE7ONqTe1W
wYE46dsmQeGTCCxd2VUawgyGatcJ6ZLYIUtu6rKrONeIi02AEviq0sN66gZtDj3a
vmDFwA/LewZvB0Pii7uJI3ZLR6ZdpeFfbmBNr+BxNUnwWVY0XllrHSfuXRb5leiN
Zq6C7ng+IvRlDUHEowk47LS5ssAhTCrlDckB4+Icuw8Pu091Uk2zgGS5YlsXaH+p
lHSsgu/3ClOsWy4+xJkEbFEw1zXOP6dLDJEoqNFR/f1Ly+OnCMUYoZ7OtH3Hz79p
uHtSmSebD+cpfT74gnBHFNT909oiHrGAZttpu0oa1L5h/ZdPwPocswMePwtYfc2W
ZAdEOxC/WN1M6l7kbENbiuYyMnRrwgX9p1oQQuMRH57o/zJs9k1jNAbQjUeBIeYh
N618j0pPCMx9EB2gsaX+nhzvMGP6zRY1r7ngh+h0nLxledbaBvMJ6dFj/abRaSwY
JVFOuE2KBr9VKqZHjVp12spv81akpOZ4JlA7o0iLOzRUZmr3KtJbm0fMNr+x9kTv
DhOEyAMKUoOtI7yAhq49br+9mfj1/U/HpM4I8a46A25Z7kBZY6MvHx2lJcLzU0ae
c4vcSg1uZkG5KGhTG1lvpBV0QYQa/QIYqF0FhPsSwSTD/HrIAVNSmD4aGIUxuxC2
M40v/V/M7FLGpG7CvEOLXlkurRCksXOgwFH1AKGC3zTEARqLPP6+N9hLsUUMKwIJ
l8XCNNXTQLt4/Gh81AzzzVXmyb+o37bOaYSVFRvbXjJIefeAdL7drUied/4NT3Gr
lF3n+1BLNayUil0T/IF09cwvZKT1mJTbtGlNmBiqjulZ+X9Q/I8nnt202OMj/1Xj
1K/dJ24nGddUmy/dQ1h7M0qQuhvBsJkzbJ1xjIgX6Kax/aQE1G1IeMjULS5ILyqF
DPjetlAws9m5d6v2KrjhxoZBa/JYy3VBxd+Lee9Q3zBg3761U7AP3sVCUHUJBNYC
dJ7EG5OsxyrXHlO3hieLW1It7aDl/wghEvfaFGYw2BZlwe4z4H4LiOkO7VnFAVNS
KvRuoijqRUifvbpu4YJ2eGylgx+Owg8jYhBgmUEiK6/fNLS+k3NuuhvkUC6SEtqT
6rN3ZxJ6sEgDN3tLA4OYS3Kr3OPWWkghrjlllsFCqkTPgMZKq1SCy3YEoZFvrlA1
Gsis7G4kSOsCnnZMQM1v4tlH7oHYbRBj8G4j6H699PcmU9wfAcJBkIcFSsrDP+ku
Mbt9S9l9RLrHKb4e0rtuGU59iOmbfcqSC8r1JNjN0MW0Bm426Lqc4Jn27y0A1xSQ
5H757pBPMAinraGbvyDwzOfFwssfsX8mpNBZH1xpyZLgVB4fwcLWo2a7S6K5dAos
GDRjVkatI5SUnbAQq4ZdSbfFcxS3lGQRh+TziKYgR4W7/R1MuW07CRsVy0Nrrk+0
8YGwFVpqAVo0V4USdFyo2Tdq7mw+A1ZgjYXQ8MjbDGQAFynmdnTsfe6Kg9Fo2wam
A5nu2tZwC1DIQ0hYe66j6spLSSJC5T5t5oGrU72t7jtOJCvNc/UE+7MGfhxHIMCw
ooUek0c8hlKh705nOuN4APdBvNh48ttS1mV//Zxy57YqaYJbt6teuBy7hYjMALdf
G1Cis2/TEd3wqHTGYelTtgjUUv8ySlLb9P9w6PdcDX5F0KbYDdkTyajPksu5C8MC
Qw8FAUP0zWw2IrzZ5raqembDsNK2igoPsncYZxLpfEdJPCj1yX2r0EQJKCjIvGB9
4rqDJt6DmCP7RPbxmGp1DwHYx5uYHGFIBkVvvatSno7x/mLCN4k91nK3WojorE99
nB2dolSPVJ/uOU33ixhOfW/oF9gMy+HCY32eWeTS5/XJNPHbfqJ/kCmSZt5Ufw2j
Q/LgRgdxZDOuT2v35akIGcA+tfBCb75JAQ7WfmFH7otr6fKHPo2ui4Ca2JeysAta
81ZU30O+b2VSB6WnFF3pjUzJn5j31dkP/aBMkT6Lb2jxcCC/cHTZl9EuEXnFuxnL
rfKTtk/XHiErajqEq/0Pgj937/ivGOo1yymhzucLXf3LPJggrRm++et1c2WwVzuY
joq/D23jNXo1nz5RjOS0pINyAPEz8I3htpjnV059Hbc6TlKMdqUU19xpoQaY5+zE
nyJuk+iSbqj26K0lInQzaeN9E6k18ixy6MK2jLFX5HjTKLg2Cd6SotpT17mqX6S2
508FXs/BNpua069hxhzVUiRCWMMnlInt7rdbvHC7jZQiuDxkKPBFi4fe3zxfY6sf
ouZZ9swgg6RlYBrJz3jYMQqMD+g/NOc6quTMb547cyPnu/9r+xwftv8VKEhUTvO8
fwsmHigEWA+ZfiSf4FmGehFNSVr3E39qjooesp7BYY9DF5M2ArDPupuRNRhbv+Im
VeWt3+bPe5Wk3bkXiU/ylTfU4sd1HwQwCuerx+DDrk+IfwlwVIrdYZoaYV2UM3ZV
od0j1b8QausO6YFyPMvFhY9PN+SXKZZMVOnaI7eijYc6ToPADxB2kOu7MsYVAhJb
PGr2jArI9gChqAA+kdpvlzfSakReKw0Ic4tWKprcF1/SfGXTz8f3mZxfIKsfKhe0
da7Dd5mAjMI0scLnheBppNaP9ezjLp7/ZkW5jxJcpleobIUuyG+K2QnTQb0GD2s7
S4VCkfqu5Rn0dmRtOIzZ5SB/xdkfqaBhSZAMYjbJruAuMKELuLdpCapzD5/8dk0W
2G48CX45J5CtybRB4Nsl9QCjCWyG6ux5kAOunIUyLDsiFoGs/FbYXngBVz8xKwZB
CX7xeHGjGq/t1z8NSXyUX3I1O6Iw5DMoxpfo2KFQTWZgIasOD3e1+46udr1s0lot
N9Nqt+MZGIiZBnaRo9bNRKlVhekRhAr2c0ABUXowDCR4e0JM6UWpmU8loh6c2nBK
UfWj5vxeHfOis6f6faLz2q5UB/LVT5lDrFfxdPXgh2G+Q9WoMnMktb6gGzafrfNG
PdHi0euwbycOWmC2uR0k30pPoLTDZsj4pBwFccMVaxbik5pjNFEVjYqaDNf9T+L2
qPEIwwxKEPQPnN4DyJxt+dJPvT9B7LAT6KmzBudVWFg1cwe94RaGfIPzvFLw73Xx
n5noKuecEluUVq315jgis7FlpqVPy+yrdKEYHxwZIUmdTSxLyfz38lQYAy8z6RMD
hWNT/TCeANdaJfA2IAVWoCblxjht3gYVywISprfyrihk2jkvwjry1+ifG+Wr3fVK
i+UzcSqJkqXd48H93HEou5hdj/ql3iKErm5IqRW+s6xj0AMi5g18YpwWX6kBCqxy
YriVoJVt0qS5e3KMZYkXy+NihgFtFdRGb5uy2nbSegnOz8viG+0u+CwydbGGwamG
FDN8RYrWQ9lOPZo+/1eb5euB/UIxfg9D+q5OwExukNUATicQtmxrONzVmq4mimAo
Jyl1cMjtfATQcZ+t2CmrZCLWvfkBhUH5vuMwUkWONC+R+LCRiJNl8rgSJgmStRyg
jSNB2rE2sK1ENj09HBdESpbmvLSC9jWBLTVbq1MSL5CvkwpGSEvT61MJIaFep2CV
kbKlP+scLrsT4PkB8hFSl8hpAHHkoZ00uZ2cTKkTfufMcBMeip1B6djNWzNd1u1i
rIOdXzZeiU+CNo3ZFfu/cPJs2YtwBaj/n6IDd9WQs5hLPF9DdBItmsOlXTXlGPF0
SusUio5WzjeImwAbPraBkeBvL4zQ43mIkEhj9pWda5sZTtKfDV1l3zn6H/kYVRt3
EC7M3sr6y6nbH1eOLnnNyoRhw93kBLx+SM1Jnyl3ZuuDSWvLgKkCQ1v4LPvX8Qo+
0HPCADbPDRy0fai2mr/toQlEzA0eQtKN6fyQ7IEKBHMuhSWudXKoWdW+2NCBbOyQ
hIy1zvqelVPZX7z2VY5tiigGE6qBtjmNYwJwomC5i1kNR18x4wzYNfmNbIAZ59dO
a0eaPKpN7V/VpkC/6nbczot1xF0ZHpQMk7m+bnUHpDXma77Sr3lkQmNE6CD4ooqW
o9judbOy+oFvbwR4bGTfD/Jk9ggAwlDR6Jg/BU2YEXXOD2yuyww4X23mSPGZlYp2
NN/TB5v7/kqRs/abuxvuJ6G0AN/K0zIUEE7Unz+xszp9fuCD9QEIWOWi0vNZLvrj
meWOWLEVWHKU53+lwzrE+Lr+ia0i3Db3KCGurT7uliz/xY7P6q8j8NZWBBq/yBx0
XKBh4mvROMBJV19t2melOkOMmIXvyKIfAuLKmMGkMRjywGFCG/nd8qGcTZs/ll9I
FY1APybzb9pZuqWvtMblBdU67fppMAf3q/Eu5LqpP/ygxCHQtw0FkvLGK87OWlia
y09F6dzmC/jDif+iEFVj7Q==
`pragma protect end_protected

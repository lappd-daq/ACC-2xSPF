// Copyright (C) 2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std
// ALTERA_TIMESTAMP:Thu Sep 13 06:32:37 PDT 2018
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
TATaVLHGOZ7yS9nRoYMuBmXlaIX/wdQJLGAMlrdKGKZq1dpS8ovhoHrbXKkQX6Gr
cudxJYoEKhM9NpjUUj2e10+gECadKpcdvHwBfgkPa2Opj0D0cK+Z8P79LmvJItIA
UKNUcBHaKFC4qwb93rFhhuaLroPl5qF1TlMlVkK9A3U=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 30832)
1a/Jbw2NMc7LBrcNwLL6g4prNfUkB58qLITYElH3cyo6AHTMWE1qKBacwAL/mgDB
RsldHHPLMQy1RdcRk+J+nDWE81C4+TWl8sKukcRr6CmyWm9/JTi2ngZFRVqwwP8M
fpJJH7jxfOhGwrezs2RbhGw2XZWolaOZIyjEzVk2YF26jDLpLKSnpK4cm2IqdMeC
dU5xeHRY3k77RRkNWpaTC+lLmVIG6/HQT0/qJS4acwRU00Nv6Y3bKjiImD+6tqjc
6g8HpcIxPn3IrzgEQarhzVzo9qXm6xE6pti58XxK8UkaqcXnNKwzCtx4OKLVAj01
Wnwo/F5/72SjOVLnco6wExKgD6YJ6YNNfZbQyek58XmutKsBVVEnk5z+n7dxYxY+
Kf2VUO3Ee9nB+vQpI4YD/ewmkHqwp8dCIB8TaMNb1O+Wp346pzgtvd068zTut8V+
kfs3Cq52ilDsIq82XZ7/HmS5P3sTz47em41/zLF20FQEZZ9/mrL1i990dk2iAkbN
/yIyLuoVhcy7WRmRN3d1hyEKbDuisLA/9O3J7NOki6mAMioPFxbpfZbVVK33aaDH
KtqiMMkIE4Uh4RCpppHr143MCE5SQ6eUoLz47vUKM6E8HZmRKyqlt4EYz859zTRX
MW9clE0jBzTRSy0Utfj7qEx4iskN0GD19WuVffAxbPrbUVwBn79anYrYtpY7NOJR
RHzhpq8jzex4CD16amY23k0PZc3/AY+f0Cp+tNwLcXS3nOht5w5ha59xryYToMdy
JZTc+f4ez8b4HmFf7bh3rRXnk2R1vTXtTGvIum13sGrsT4wzi6YqN2Z2kHbPRc8y
/DElkY6PGs/REs5bRPh7Y+o92C2zE+O0D5IwmhdHmQ1yWhCdyBRYy3gCXpQVQ8xt
P8jF6hltvhzyQyhENozE7rrNo6a0OkOmocqBmWs0qGLkW/mGwBuOSEJ947YXC98v
99u5hCDomuFvsNyIXsRPhTbC2WxphEKhnbrV688vmXsELBppsiaKiAlOfanzwgBn
85ZZJNcB+xOovwUpCU0rV9Nox8+RcdeDr2hxUiLbyP2V/Bv3B/QJk7HSJkZPQWMZ
5eZS7vBPDKqBT7n2yfR94BffIK1kYTCQEtjFsSFOqQ3PMAsL1vj1ms6O5TCAVHms
A6TjnHfoE8NXXVC/HdUZgK7dtywjS91E6lVqZr3kTVdAPOTy0eDQH1jy0QegCYeM
PKBsXX8H+LI9jBvaJJ2ALFBgebdpDLYsK7rBJZ+WkRv5wVtK+HagHiaNdX1auKGR
QUcRdng5psCv8WHYJnJ8J7eYKrvTWxId30xaYyCP0DN7c3zHjGy2oE/AcztzTyHo
E01/nWR4u9SG+o9NA9UJS12tdpUvtF/9GDOLmFdKtCgJ6+xNVs/3Z+ENXGAZO9WO
IX9dAMTHNE49Isn8xj3/mkRG4p1hODX6CsvMA49SZ1QfBu5ryS0+Y5vknphoAPSS
cFxl2ZsBA+Uns2JdeAXjQOqWBriSXKq8OPbZmocq6u0fuiD2rEPVcROmKtvDDkWO
jd3si4qQXNeXT2ApzWqbnmfyk2Kh3YFjcC5jiCBMITsa1UNH0ewDcjd8AbyNvuS7
1e0qBGqxrL413UV1F1lhSsXy/1hGyI0WJ9Rz3Keh61Lt5AxyKG1eEPpfpdp0sQyQ
fV6od319QP4s/MiwMvxOPp6dJu2JFo2R9bKG5moiTs2q+MwrClX2o5v4DrUD2Rnx
Dm9bEbW3htezChZT5PopDpsKgiwwtsMtIBeNmmB3b3qlwS5Vo9JaRXcPYN6laJhc
gG91LaEUKc67ZJevqXIG7JTd5XgTc3EaxyCg/16ANNfpd4+IAqbh+QVehUXfvz4t
6smPB4K0GyI/R53525jyuUYyzDHR1wSbVLbKV/inuClIW3PzXzh+xJt3iKcHVfOU
OyvwrkSTt4M+p6Fz0LEBYej/r9Mjr32BTELYxV9yYjipp2DfWcqy/kp9U54dSuRQ
pcAMSmEAvUfWrkQht5Ka1E14m/7AmNOHXJ9ndjiNCEG+K3h0fuy813ke3PLDj+eW
OFydByQdxXmmz+UVg5sUxwre2w5NRwuY1XalFeeIpLS5z9yqcXumjgm38ATgH384
RtpEX1ScVpIPifG017iB5m6x3/jzSTkXGYOQH5ir5/pjan1EjGLPmIr51ialgQjG
z8iudPF8t+HS/bkQxxe62FsUAKlJQXGVJphP3VooVUhPCcXdarXM3pJQxX8V4Vjc
RfCgQC6fUtM/7veCMppmnJI2krkgvr/NxJhpr6ujZVcsaQM9OjfEUDmhiaA4COKb
bGLbcaOQA36NFTuNzXDg0bVFji8DermK2ET73lr+jOiYxoZZ31XNf2X/z+Uq8oXO
KsCqyMmNhtyDwdsRDSFXLU89aVjfr07w3LV7zY1fAA+YuRoFJ9OnKIwmgoDJMrsb
Jv3tJrucvTd7SIkpCNIySXHKbNi6vAE3u1PPYHHotzCEpmDTXbzF5vWg/UJfhVaX
BcKsxIkRYxMeGOzftInKmZmAu9pHWy9PT1dYzrau0tNvmA5RlZS6tanbacMZKHy1
a2B6OucsRp/DvFxB2b/dQiVbchQTiB1ttGtkiTwb+PVY4/AZtEXPUfN46aajus8P
PHvaZZdLDL9ktEA1Ra7ziUCojd16h+LDIMPv1KYoIqDIOeGa79+eHwaZ4lhJekcw
q91j8O+4EY+Dp4JGb2Gi283gly9Kp+Jncv/wIs1ToTJyNvrVc+/4LpZ9aq40MkdX
4vSODvZeOfhbvRnHri3HO4Nyu130hO7ml08aKrc6ggo7/wZzL0tAL7QMmTL95aDQ
mVenv4UzaA2teiKr9Qlvl13buJgN2GkO0pPDtGnvMbzdSFsI08K3oXTtIfvFliNS
RH/4bzhLZgV8LZpHh8YkoHhC/NiKF1OZTYnYCpJSGO1Eov0HPGuhIQ/O9f5i4Q0t
a1s7qNqVjjWuy9BXQH3M39qypGBWch2s5aYyhsV+IJqcUbDTMepyhRgwWrMkowD0
vJJO0SBd4NEo67nM7AslHjUOHohpxaPN9gGkta1xBJiq4FcKRK65CpBaFmvGQdxK
R6YSgwxplmFlwYB/rg/gUNhb+OPFrrWmKChn0/5b1Gr4U3zxFj3m0pIykqWOdI15
N/0EIE0ip/CXGYz/2JFGq+W6ougiBvyIf/7YJfizKSgW2pV94yc9IhnyBgvSGeaY
tD4RuGejBaZ0yM5rGUcfvy30I2F7vUScL/S5r244GZs0+R+24ZxjYEEwJ7ATrWXD
OIIiJGbULVdPFQcnBVVNQXzQR92crsCDwxpMJ9z9ec0bWx0uVCRXSFBqDJ50qSHs
ERNr1Z7hmBh72twizHKAflpdyz7FZuWd8dhpc/ZHyCge4nDw3Fx1XS55fqywYsvE
MxGNU6DaWIej/JzNy2nPrYfBnwjtOMmFiSkbbWlspbI8jSeXQ73MgYvazbLI5dkU
FqoHBuk1ZjzCO/2MrAFqleNz7pCFNZiIGx0UW8U7+OZc+Z2Hf1o6WsNFPozTuxq5
Y2ZIri4xT+rnUidjHcVhHu22893g+tz+6qPA76hAkiJoUFHhMw/sb2qibqhcO4U0
uImxuVCrCb4jX4GNJOJp47NCGhChFSm70Cru/MDVS5sM2l7kur72zEdkD+hZ2VX+
rKBWgEe32wMfbVFrjF4ogU1WFDjhg5S9w3h/o7LdkVdm0uKdQQaiQhDnpEpVUj+s
IApgW05HVXFkMq6EQigBDguRY4JSIDmBTIGfIYKTokyfhAUaiCDlCch4hTFxQ1wm
P5DbrtMqYnGefGTg5ZyRUFsy3Sjm6H4ybpqljTm8r2kWRMkxV9hZ20YbfhNGtQgW
z07nMUOGaWZs5ekle2seOyNHeMOM62eDw837CwYOv/PFKbmczNagJe6Vbm9Rpp8e
w18tmhbo58Bw+cmZEDyB77djucX5E5ihWoAb4zfNr7EKlBFtlYIrqoHHghNNglPJ
EKC0sLHQ6GORJt7HxaVKzd4LPjYCduA9mrwStfH30JiVOLjjQsqz2FrgqkgC7hSB
oeAsOBOSf2mAfoQslRZ6HXxqhZmJHj0Qd0nilO9INe4NFoQr7MkRdisqqeVMLxIm
FRNzQ6usq2jHSU3Uxt96AVPHbvuJiiPA7Uat1V/wNzzrSTMlw67yrWiL7CleG2WE
pSxgNssC6pUkhePHOFQS391rkjgAdn/Oedr0OOjsAOpugOMQdds8LLG20dZ2S310
D9ec18xOSqCHp/ULnpav6tOwuqVd4sXKUn2Y+m+AxJrMWKZIHTKa7ILhXelcIpmP
AGz/oYFVQlQccDTk+w+6AXa5zrhuFSIzd2hIwj2IyU3HOVTc+ysvKv2LRjjqtOYd
wgnKoDDTSRCL2WtwoEovbNpP+TGCMFAphNoXGpTl4qwMYIVujHNP1efTMJqT5Gyf
ZCexQVxisg5jLGZJdc3wg38Z7uKi1MIX9AE63xy272gRqwQCEKx1steGKX5XV+u0
8VRPaM05G1OuOP9HhplK3+cX0Iuo3D+AGiRLJhhAtCwJS4eiB1CqxomcI9d8BkyJ
A0mp433Ba/cLzt1hCf7sUSOb4A6eBZakZKKETf8A31Gt08waJJgFf3wKu4s6kzLj
3uPaUQdWchASBrU/QmdRFfJSmumGAnRt5ffxBb4Ez1lVcrJTIVO8LuQ5dvZHBYu5
kpF5z8RcIW2WAiNcTq7NOc7qfqdCSdBGc8VCtfSw7T0b8fm+0vIqtHyH88aD9vTJ
fw1RU5ifraE4rL7TCtNWTGQRet1GdyPT3nV5yCHSYkG3pUpftnBC0CJKUCHvWiDT
dZbMvDNIkQViV60SbXBN7vcqoRFg/XNh8617Sm7JhPfzl7V1sWS40zzKh+TBmfqi
2eV5MVYveyEAFmMVkaa5gG7r6Qmgpb2lEAkH7laAubAsGmu01iCDY1LKnzCXyBwR
/fRyTCX7pDG1p88iWE8TnzIPzRubNZhiTjsTtVX2W5jrefZrVKjKixAoaeAjwtTr
Yq+La/Dfmay3bmCybxrTLYwVLE9/2y4xdcHaP7qUXbPsm5WKt4vhELPsSndMISj0
6/U3rUpBIoMkQjZKAGD2yBvw3BvYUI+l302XRZGDEE5Az0gNzuuVPen3ghdercud
TeqoaeUlPQaKemt4O5KlhI1aclBVkzr3uBceHF8t3lTRdqdnHZ7wWP/pAXHYpB5P
fl2wIxKQwXywqblD+eZkqwbzZlMFYQ78RYmdxRan5X7zBZz0qpeTsUZOgZwdZMBo
2Sxo3IGypgDv/gsIchFtFp++6VGtiExSaw7TWfMSewO1G43CPIegrcNASUJzcjWx
yeroxXdfiN6QVpKM4OUfXolALP1DRdtFkOj6AwiQJAjnAeJQYYprV/UYJW05ZiPq
bI1d77x3UjtejHEGovBBc/3mU3MpyNIwsWOGLO+GRh7whpvVS9X5wsIfIU3vK/RR
Jo9MlLv/Og71CNfZLHdhoZ9SPW3DM3W0Mv9QtDk3dXeydheX3OeuTXKbMMH3b7hK
fvnq+F6pylmtdlv7dO75hiO63jX+b+IdQ7fmDLjYeaIQZqV3zvRQFES4br4fJNmq
DVUHStRU9Ku//3rmTCfPmaasEyuRAEri79QH18kWgP0MoevljjCb9M/PcBHLe4AH
fOGv8SUk0jImJsrowNDGgSNfkjM4hvM9d7D+5gr4JLwTTToiJgMUbLLku395USGq
Gz1uiTW97c4EWesl5Co4x0cL/HrtT4zGmgbXLBx+AjvDPUD5g0yrSfUcH55G6/dy
FZyIvebDSA4k5fqf/vBB6eFuIoLWEFIHpv3v3Sxj2pFQuMEm+1T5tGYMOVLb9BSD
KkLwCJWLKBp+MbulEGcYhkKz0jW0DCNCU/90PIAfI7Obd61C69g6rAGCZYHRKpIb
BGPtW9wTSKjBmAMq3dT28AELa+iZWXO6D+Ze3X+bwtBF09yEJoKZUXVI+i7eq+PO
Apl2xMJ9lMiviVPvdnGD/2lutEtYPsImLqdBikweOje8sfsf6ANNTxlBumIZnpf8
TKNXWk/4esGOW9gnB+n93R4IDBtoJ/FHTXhFkpLwUnIB50+DDbrUDt2R8hhpszsC
dXBDlaAIKfj+6rIxyyNRX21FbFMUsS5WMtXASHdiA61XaXn7zfehFtHCAqfSVysr
6lVIdkkxRZqXO0eYwJLNLTD6rM4bq1+rrx0BILboa1kILJlfhxP0aFvAJoTsCWEu
kCRjZDbCvZ5W1wYG+fxJVqKtFjXQL80xivDnB/0hh4pEhd6IbUAOL5X/o8l+qrxd
jlnmgmmxIPm0Ch1pxKYI3JGjEQ8HNj7SxVS+5svCEhligzs2u7ED/I8Smezd6yKK
FVridPLJgrExbAH4LALB3o1daqojcG16APNq64MgyRLM+AeqqrOSvc/TcqNjKh0D
2Uln5HXTQ8MQ6rY+zyI+BxB8eNpzQFkf3XZEFNJmcdQJDdVXB5We/qNnVB0mpw7W
EVwnrey9OxLRKDeL1+e4DJeS09FZJpUTtPES7Wl/at/cdT+lnYL3KzLMdYnmGpIb
JJrglL/9cMap3f2qivWsJsxDfsQOl6MvZjr8BMT5JHi1QVZSlXIfIvaKW79csKoG
Gbkc7UUxJU1rVCpWvrr5gaa8z+sttE06Ww8H8mQfmVdrQrcPIkIMwAxDMnI4iDqk
bNQtCfO+YqSasEsG1QXqon+R5d9OpBhue+d3jWUWx9cbBVErhLgoJRDwHfQc3yma
xVjfnCTBmC2xALpJfLMgoFGXKseI/aNxMAlG2nGSOrrB4jv4pbq57esVwV/V49Da
5ImGFFbotJg2ILMdOAtyTJlggzneE03idGCLfYV/8eayTOuIG7YpfBF8cbG/gF6X
3vleBGtoARo2DZk0JNqZbiYPeclarKy+qS+k/MSRwQqHSmfAthjogfH/fGYegtFq
l15j9aRH+Ey+V0lDzcJnp75ER1q8HhfbO/iIxKSgzQCJDLUeAvMX2kZ0jwQW3RJc
rBfp7Ax5sEfzJH9MrAa3GseBhyp+iPn+ibOU51A1L/hoLf0NvicKx1JpMYDb19MC
bCMXXOlZYxTdTOAQ263eLzN9GE+RYuHRlHHtBganwfb4lrSgJOoC93t+3ftDQvPI
YLYBJbNZKCn3V6CZVnJgANWWwKbS26hvWWnygm53Y+7N1IesGTOO66V1pkhOxVvT
HDI6NDLGUc4Zd4IjUbenmxBagY2jFURfUfJbm82j/hHhsufH9uJAM/w0kIBtOXuC
Yj6TQz/JZDg+sO4OU10iSlBnsW0a4b682fk4DZbr1GQ+4AKTm3ZM9dZywgJFF6rR
pdLXch7H3ZQPQ/de40MVL8q2DGwmYM1rbfNeucsZOA+roXFFJLY6opuFzZuncG/Y
wxBwVpzW/FwMUqI6Z4BCC+QVwh+JGDDdRWMBttGXIZoGLxcPzKcUu3KE7RNLeto5
dT/KLuhzgPGwR66K1omKHWp51zzMSejLo7C9dZq8iZ4Anp1IR/s/vMWZOj2W+F80
zPQ9cx0/vFUrwzHXQgb+KpqSmleB6+uBtYog6+YF1AHt7tfExQvvcFGvAjEIj4ap
UVR0PuV0KxCQMV8y9odZgj2Bnyg7ncheLQk78fEDbjTzk2F6n3uVpD29/UpGz+7X
1BwxIm+Cmp/HKET7PzKqjBH4jr0cTWauiC4YJfnJLD6SxAD4vO8mrCGWojKiFhwL
0IPwMEDadJU/DwEnvlZOHjqXiAN8B7N82ByBaSuzr97QzJUsAdSELiTVbT1+t0zG
gyOBOk4cjnVUM75YGqHhUmFVB3Hmby/Pvrt+xbzdemmZ+jZ7VLUq8O+RkpR1rFz4
/n2zt4UFeKXfeNUrYWTzE2tCu7cpBBNDFHcpCBiuTfcYrGparkLtiDxnM3u0VIGi
Liz4Qu6C4dHxViA8r9JLjzznr4c3HafwtLuDF9JLF46UY0sZ8HjgFsHcdPbs0eL8
jsa+zb3b6PP0Tz/3Fw0eSb0Uz1Ac36/pu9L0q7ZMvPLmAfhyI3w3sFxEWWNDNII8
NSr0N+qA3uh/Z2uHnGI2WmxacCLyXfaVZRNEUZHyk2nKLNYIJPCzgrlmFsTc3p1d
7U2FMI2sPKIM+b18JRbaHWjo2RCnKgEdX8rXEpkWIjeAw8y4M28PMfQbXlG0wNrY
OAH4GFM4xyrmCdrm+2nT2tD+G5ijJDVD29rskrZ4fQttSmABGfgl/V67yUDJcLMi
3AV2kZtmlFJ8A/Zj/zpCVBMSr5keNQj7G3tPlaaIrLlszPGRb5iiI/oCDmOzeUss
2/6nmE0hiKs+BPUxBk37VwO+IGocoiy1EPXiK5g88yen7fTZAtrqx9BlTen3L4pe
7RAjLx+oH/zznGXIaypMhekxROa4ojpQ4xcQsQr+aBrrBmpUlyTfo3YFDdj5E2IC
uFu/GNq6ozE5KnzIcLBgbCKX3YbaUeP5lP/xSJu9TkQ1Mol9vZR0S20suUJuYY1y
4//eZM+AFSIE7IVW9u6Y10vZMYTNxAecwuLIHudUbnnfyuRQ71EU7GIwZiC0o6jY
DOBxfC/VOLTpko5fEx9cOZyrnlkjjEiPmBGcZ/3F3Gw7KPNBsQDJCqmYEdSMCqNq
0lIqEl4eKcj45IfKdxOqI634CLXB7b17D6i5PearsEle8LuGG4unpU4kZAP/wQ3F
fUzzLWgP5lQ6lb96C/YA1cQ6+jI4DmAzE5UuJkDuv3iknzHdmpG5Gn+OwXUJj1pT
RYqooHUXNT4e9KSVBFiOiQvh6AArxBCLIt/tFm0shsSr2BiKYyAFEOOnNUOYTf8z
ct1KN5YPyBvKPxv7hLMLM+MjJXp3DJjzK/o2yhqKejkyLCJ5Bi9DL1Vdf0n1hIpX
eAws0l+fi0J1Ubr/dJxBeeOzz0tsesTFcSswp7X2UXhiRlULiO99/TOfvPvSVYWe
2y8kJwWpHcEyvaAkNRw1Thf8BgTW0K1lY7euZYxXpUA5C9/Kzo/5dy+lzUN/SfTS
Fosr3om6GgjmxSW5c3X6E1r2/wPoacsa72uw5PsVy96czMJS2d8leo5mRx/nEO6n
LzfTtgKbXJpp16muOxnH6PrSXeKgQa5C70BXsyd8k9/kLzuJzUh9B6OrlTDwJ6Eh
KaeugkMItK/kfbF4O1hHrz1YxszG/zIEMVHeLejn3+cwbPQFJypgyNIlrRMfAJ5o
7zHnsD4H0L63fRiuF6mZF3jnqlVn/XPyA7wj9PtsVuQvm7vq/BRwCpxHLdAvHgkn
Ib6ppfqkmiNqpI4kuy5+VgMxLQTclxQXNDGvJpafZDGoqw/aGzE07usevHh+olYk
Q0I9utE2wzjh1GdIcFwMJdg2SK9UvKzn3ipBXh6Q/VnggzZgvgPWoybeHXfUeSxV
fUb9xlQb6h3P4VSairvLyW8ZrPgRXdD9w85nPk7riOrydYjHB+ky6AiLw8V2qlLY
fIrn0ftasE9gQDRzDbe50Eprl6JugoCOby+UPNOgATxnbh3DL/svi7bx/O2aNaiR
r5McZWMJTiOKJfQRxDqrIJcgCzaIPootC2WkZJMnJ/clpAK8TifU9Go0MhJvGP+3
TkrFWXdMoG19s3ZkgLV7jnh1DV8G3WEwalUwdUrJ1UaP7QKVcSASMsBpSkxuOJq7
Xwbj8ie/picCWDkxpm8H5FrLMqKRH2hBuPHAixUOwwkzCOdmFr3XudMtaYSFeUUq
c/tzKxtVdJlXEFDVgV9PMDnSpZH8uGwU8gusbRNa5qLa6d1UI3seIXh7iTDdqgas
xVcb0SNJPzFQ2wbFaefveipUscW/+fhTLWXK14Hdgw15yQRLJ7M40old108FfMPU
RTXVnN1axZ4oJX4xCBHCAH8SFWlorhdr05u1YteyB62zMWeyKgGcSGsVainrQMWN
WDnjDT6vv0WG9BW3in56okhMPCk4Fc/gRM/95RW0WICl5gP93GNCklcZgsuuH4OM
0PqxbmNyo/tuIciz2M/8oxpJjnGXbRgd0YAO2K6Xq+/MTE7BL1GTpePHPVjfalIc
+OQLyQo5nXV8ZptHSKLwR1MofZo/9jHPbIzwHjlOyv5Zbr/pFnYkSwqW6OtUFPll
HbLN7mqWbfzNI/nssZPwy7t1cH0JA9+Yi0VjZOrDra8IhMQUgBYVOfxSVYhu9Js7
5GQyKrb6Ca5iXj6MfVSURssl5CjnB9FoZ72aViB7mHjtEfYH8YjgeAOmkDTiJx6c
/JB0jKjwfriLytTOquoYtE9NWsEv61LGQ+ZDefaw+pkr8aR0urt+vmJYc4Pij9Ey
w39GZ5wlbLf+RlRKJ42G3uStvwDaiwiiHu6qud69oz92kBhKA7DlGE4WoyYKNWvN
kcIxILsrj2QGp3l4G8fQ5WvLfDkNrpkWIyrp9xWs7S4vff/curVzgCM+rDAUyijg
9kcMcnW/neUgWbD+q6RynqDSQCQrjIfe0h+AFwvFUv27Iejy+ZeTsz7y9m77P94l
Uj9wKXGnChZ33D5BaM3yFXtM3u15kJfvIhVtHqcHj7xx2/LmrZnI/+XmMzVFNgcT
6CAVyB5jO0q0TSId4SCUEbe7HkOsWmcsq8mmBZGyBZdfmvDzKauPAzUsmVdkaCGp
Q/jKYMdj41kcEr6RMWR5M+NtH3pe5mmq8Xme32e58oSnCQFN1LHjmd8V/GiQHn2h
8OyAHpoHHGSKQSXHrhroy2Kyn6PiuNyb+g/f2RFmViVJiVCz2+K8uzsi0TKklWCS
DqrD2eevMvk5h2yuyCu2k4TGkyhfI7LxyBjpwRM251ZOoI5AZxBAXc4Uc6hf7IEY
IaIqbsZFjE2V7nHZyjBnqQmY66IqbDJdEooFu3/9f7JTWUK8QYp7Deod8zzMpqJo
HB+UKfDeN2+CPNQnd+XV/2NUNc0+WJht0BO+tN2CRiWXOk49Y1PnBkWOpMBYSg8d
zt8UnCPmm9CW5NXiSLj16PW5b1am39CWSm2US/TMq3GWI3uIcyq1sopUC2AVI7Pa
SUKQvM7YQrdAQoG8O3thB8fiLBZyH7kSWZLz6QRY743HPSJZWLdpUROM3EgARNtz
mGqCXVYZAYLsx0fnhn9ySZeRwiUVgzcMbo3c80Jyq97dtdC/ThLF87QYJTr5hDn7
IdLTQWOU1wQEL6nGwrU9n84iKrJQ/lHKmdXVOlD9Fs870J0BVIvQaMp8mL5mv16u
uJ8ZQJlitgCSteQdhkma0n1gqprgF75GClGug1c5gKVD5wK9sss5j3V9B6USzqBu
H81PdSXo5620YjGjveG1wRfMhe9orQQGNHmVoz7VDSm32pQdxjfzljMfFe5Ksqtf
l8+YLy6sOzdMPkIIrNqf5elDAC0Fw+hUkrW0EnkK4qMLrQlXa/BShwjI8rY71HkI
Pifn1EWHuNCDLn+MSYun7Bl+LF3G8MFucm6sDGBVe/76O4g6NNB1CRh3M22/ZWor
FX5ekXQfyewMB0iIgbAHLAcQV3LthNVvznEBtJx5/8ZH3GIWmgBBPOaH7D1olzcg
ncZzlmxUbRlQWlBK3HSHwfLqNMsGQFzkZWJpUOTvBFGVVn9JOl7bpeg1wUkFtH4K
iv/Oxmyk7V2+bcHGkbeJQI2LEFe1b0zhTHaLJTABoNbJZQH4Mmr25Hjv+AGE17Tc
9ELQ0lHTnuTjBhMxA7NlprcWzLLdoVvKXCNpzToizGI8t3pTUYf9JaBhdMrM2WoR
bC0Xxq6ZMOpaT+KFW5NIdiDtgVSSk8KZyJXpkU2sKDshLVJbpVXtnWPwilyjlZu0
sr4cbDwvV2ZCfR8UbOuSW2JUdZ+KiYSYsIWodViJUpe0C/RCn4praS554K7KhSp9
+xO8WiW8k6GrDtQtPEdZXVeJ9r8PMmMIPQdfBsdCdGzk0qEklb+H6J6ospJVpCs/
RSGg5IA1jAIynX7X0vIkXCphxQnJL6DpJfmzndJR1+l0Grp7ii25Zs3+dDyDUmd/
64aD9MHCaPz58dI5WkIa2/+nISROlh8nG97tukxEDTTRVYBIxmwvIRND7vNkdZn2
71PB4wf7P9dhxLPSENG7czrehGFNQt5+1KDDN7iXBPcjSNQ5y96IhTpxB1+uZ2xl
/9flkaEM7qNZxBpUnCVKyaVONPgFGasONZW7+n3/1MFpVvvidCDgVdqWagsGwPr3
/I+Epu+FQjAzzzICSy363qQZlzUL+NU/J0Oruwhwbza/YWd5bWVWXvnXvq0BD4/z
hO/qwOLkssiiNkophUcrj3ngEXluFO56o3jri9nfuP9r9hNy8DDqe4NiIG5Fb7qZ
Mt0MpudEE5eO3GeTuVaHyFJYJUzzxQekSWQJNegVHo4l13TIdHoW2ktxhNLCsVYT
CKKiIp88979nLvKoQPeurg/ueDICoxkPZekGxuAfphcGqe22oRtqEpyUrjeevULC
O5VXF9WoQFqMfsPk+QKJS98f2xvvunbbD4kdUTi4mCLL6jnTGfd10WAMyJAYwHcm
FdN6GetyX/QIl61l5anNw/EF9dlPg7a7NOPWymP8Ox5efYPjT5M9D4LQn2MsPcFr
XvzwizJwzALOcyEeAGrkEgwuK00hfwik4pHjXjHAAg4QLjH4aNqES+zYzQIKAW2A
Ka8UY/OFF5/yTwwoNOsgQIdh3uytBx7oy638zW4oQpDjiHxdtQHGcNbB6hSZ8CvU
GuwZmmDY/tVKH4NTWzrMTj6kP7lPGChZ7nkW8wBPlBEJy56kTjE01UUatlRABV/4
8mAb9ZkOoowo5JSwUUsiBzCYFaWqudGVf6trFgrM4dgAXIiMKbzlMacQxLHUsQAO
bjMunKSTQVlbPxnUP+dmd8vaFq12MnXCWMoV6OcwY4orHlrKJR0UHSy5hyNf61qp
yEbikaGQmhkbX24Ia/513+7dV7Y1lpVYNYBTVoGSRZ0Nafb0RpAZP1UpaQh4yY58
XbRGbAlLhWqqXFQul6W3MbKY8dOyhe6Q0EL4bIeGiuhb22ZwE2qtX/Qzoq8B8PtZ
yhMdiU7yP4oj1tEgcUOu630m/Pj2szf5Hv8IsaNTwbTd8WSsaqachximu1kvj8zE
hQoNMaIQBMENeKFywORIs4CVUPJGCG+Wnzrpzt4hR9FuJeVqXsKYmiSMKUzQAPeu
4wNhJgo5vwgcp+BHNO2id7WSRlHtfzR1Rqpln2k/xm//fB4QrY5ztl+kuE5Q36GL
PoX9NLoLjR3ubeia58f3NlNg1mg8RIjqJ9iYp15PdgILIbLJ21V9xM9+vhDHsIKf
69nj8Y37E3n+lOiUEEIUWpYO88KCzfBhjSVKSRj3fEyWpn1vYJ7gpmBvbMNKv8lH
VfDnvk5OmlsIL9leiwyeCjgPeuF2RQqtgOmrfsBKorYBK31gHxR4MHCWpbdAkJTK
bqKfoI0y+//6JHGWHWzNsYygE00mDW4/PEUVCA23arhymFgpuwq56CwNyD73iuqP
tgI+h4042E3uqRsGj+LRgUT2OaCu+d3dFUNnx+uL5O4ri+NjwSmvlAAIm6CaKDss
OXV+eH1jG8o7M80kilxsc0DDYoxlVeV993FTnYOwZK0rrUac8OBEg2Kre5u0rTQe
O/41EuwufG5Qe0RNRonrHbJY2pb2/E3Z4xksjFxrdyejC9CqjKAJmhsKgpDLP0cj
v18SBOq7WKZTj/ectp23abqVjTCFn6RXTt4AAWP5fowiP53KZACPKQTXffsDg2W1
dpkvY/zNZcnf6psTxLx6Gop1B+RpW/n77iEGVyh/+twPtau9SSXQoCRgV2xyFrq2
YFOJpWrSjJAtyMWN87mDkGvpaYhWRmYCNoh3NwSbVbLVvDlORy2cdgp26tJ/hCEG
0w3ieZe/hEW4z4r6vIowxW/7cIa+gbmwYi5819dVj3liYz85IARpCbJWxWO5D/Sl
FtsilhwL4fKbUSeU6ET7oG4n6G1QLCcCcqWogCsYeVwGhGRr0ubUfw1NkXR01WFV
3ovbojSKTLfx3npSWM4kBdQUNIV2nCMCcl3s9uL5AUFysZXFl5CxHd/trObu+hGH
oIK0ThTWdOm3q/5ni9yVa80ly+hXJF5C7oNnoJ7NJLc+M0BVaRmSeAnwvFVglyR/
DRWx51UC2aPa2tIEpDnQzRAluStrK3lKuxxcvsHpF01L6UiddstvWTfstDlK3A1Z
iQUJqYzfkaFc875NA3g9j3LPhigFHTjLQ2wOroxOkRW761Z09keF3KjVsd4bQc89
o7ytHJmLR73xlM8HnW/CoN7eO/iqYNoOp+1GC5bVv/OuHPWM1AXKw2LKvL0bqrzf
NmCay4uv9/D6UHZR83wYZPSDQ5kT8G2eZQdLhFZbxXh0kocjltbxj2X8RISNayZX
pN528jl19jXwoRtO9OyJDahm5DIJK8qs/Fzb8+TsHdjU2E/iuz30utAq0tFXvwCb
IdzKG+xssliVmUL7wLH4sDdjTjzyvYio508icNbblf6fJv6PeyR2rbfWYg5+t8ha
VZvupp1K9qGdFleztLgAUN6QN3ROBM2kk51fmI7Qomz4Uj43c5Y/7PkLguBYkd4D
7OEi5QWYxZNVBJbE/KnNxuZlKRny4jD8+8391UoiKfn62end4WW2hVrljwLZHqsX
79fqD+/ok7gfexDJh4cU5WMxaIHUzSZ2tLBRreV1cKsRXbzxZouvGud7OERKOUmA
UQ6s1GxznVhGNTZMQDejOSszWRtoZu/2vgT7AC74jChPGZ2hG7/vutpYxSTTocsQ
LIhaRA12deEcR8zfyGu41Ce+jlEOvg4f0t+utNpWiMlz6TAr54X3doItSsLfksqK
Fv2/O4lr0yRcDFQCBCUxYhLzDgxbhqy+o4BFlsKBUft9hNZcYzWlKYENsop331tB
GLqabV0L5GotfX/7ZXuRYwkOUIxcKusski1FZTZTMSVZL43jc/BdJP+KgYYwL5rN
lOyR3+AGUWBs6tkGoOO3/91HbmKjkP08KgiWTBsmYyIcoLWiNwkowXFowcpCxr2w
yCnyLpuS16fXIg/BTwfYkR2iftjd38nwgVnWpBXgx68pDGOGPfIl0beQIE9colRv
aOBmYzSukLcwW7rbI91Fq/lx3LToQLg3kvmMAHxJ+dY9st6TwEVqheXGs3T6WOL+
x5us0WDtAb6oebzS78CLaXjofiOFrX/gzySbt0BTIakQj7sflg2csM8QxXa6f/j1
ALCUJH5zxUBtd42vcUtlQ9XJ+Era8psIexmM9sedDRyp9fAsytmKhJQfE8gAGXy+
v8YOS2qEK+hnMH42XIrXXcxDxFl/UcARdUfC8WzyvgMGaosUozEAH6njZwScNKpP
d3/y3wUfqk/5ObwO/+NF2L8o9tCL6icrHHLN/yTbS0m1JUippfjaos0BZK1sKHdJ
C5s/lM8wFvDng7xcs+MBijQnMfm4MsS9k+BnD96SbyOPGGY+m5NzkCMKTFTvYe8p
IlJpQNa+dsENPasEzViKe8fETNVI79ytMOtfWT1a7drmCuiqi0j+19kg9UJ5U5GS
8UQ+xhXmGq61RZw8s4FzfWk2zsRWLyr3HxG4SfSVLR9JWLiZPkUagTw35gI9a6jr
X7CVLAhcOaq2cVtoNAhZYo/QF4tH5gE05KzCHnZoEsU8tDvOhjQ/hFva3hwKhmrX
tzZgBHyffidX7reoeaUy8zJ3ot14q7DPKUmpTFG2x2A6bubOIGQqm4jr6tUU3a+E
9i8/l5J9hmuxfAzL9Y2s620pC5RuzZZ9MzdKMHdUANTl+OU7MPeFlCNad4NQwQBv
+UExTIQWuLP0yFL43LVC1FBte/wXTCCj3bmhTo5vpKq3BbURZUKYicSaIz1dPFbM
Nrf7jGMsDOrJljdroa8NZjJaRauiRTZGmvoWDqzP5pd7949aY1oV+oTWbIvqj2Ol
vY1UrZbNX0q7A22+OgVEi0j59kzr4KzBgyyeMP2/CsHq8BCMwrLiPbSLaQmkt9xr
eMGyc8YJZWUSivrTsiRx9BfL76bfaZ3K6pmaSuvkcjFJD2BkfgrcGb31DdW3yqh4
FEP0whj9a7CsWyBcEbAhuqwVAPYtEUW3fUp4x2afJaO0CA4S1xakSc7N0sZa3qqI
P7l3YqPY/EOZz6FuirRjT4v9q/qfW3hHjECZBTrQeycv8+zu3fkxBAcVEP49+6eb
V+CQkGzvZjpyHnH/h0J8uIeR4eGlNBELIJbezT9XsszNiZWQDjYTyiQlY7vCrNAT
Wo5P6Ou306AMjoNav7+bGZYUnm+YEf0tZTtm+HUZV3rdQuPZHPrJL/sKNva0ExI0
uuRJ3tpD/9VVImX6jN/f45W2zIKow4cG9V9nBvBN9X0p2GMI4OQ9ncYMZA4Eug37
nbq1B1YIiKjOW56ehZyT10lqzNg5EuXuJxdKiM/U3UIuC7KDH1WuJkz0Z1HQlTLb
u5l33eWhdTCyyfcJUusChlD9DZJlOI9UI7beouyuvHgxQpvNqxGPvs8d1jZ8gaMQ
tzUL8uW4n0AbQvamWZ9jdaeYsFK9WFRfQSTJsKNZ0e7sEgY9aNnkNSTAhwTjpGZp
HkpDRmhfjyv0WwrNqwW8NH/f/Nn/02GA9RJd+WTNls5vOmPjMeoqVcZbvBqk+RZf
iWWNLRom6psG1pLQSON95JnEnDtIcyQS1SlaRFH4KgqcjMuZZL75wdB/KeQKp+be
Fkg3yswIHtVUO2azwresPQyKYiDdkBicoxYFEdR/AZMCg0UyCZiiYWtGNmFAzKvV
PzZghLCkCfyLIUdzsP0umMU1Rf6fmJ7Mk/6oHL0fT2c2YNCDyZQWt02Tg461o/dK
Z+uGN7WxDx5Ff/9h8mlo6VGQi123+neoYAN5cyP8+SMfsz/EwT89lG9RN2aatVDx
hPFiA5LSkI3FwXuEpsgG5h6PVE6H+Cj8y1XpHaOHfs+aQupqcOhzwjjqB4ekHVa7
otIM+kcYPZNM/JO8wIuDOe2ulwKkXm5LRRuCuVTSaDO2uAJXN0ZAwxpmcF9Xmd1D
bBAB2rPBewZCaWoiDwOwCaV5n4HrC25kRX+Aq2dxY6vS2acJmorhMneGdv1Ib50U
+TFZZYoywEoWHYV9uAWbPKiQ3HWW7F8ShPi8qgoTHMb4B/hv2grk3CgmxjrEI8a+
gZmr8pFafV/otFHr6dlnzW0/BtV1HoorHXII6WnQ1UBTFOzMGJnl9SHEQMQj2rmt
LD1B6klXvJwX4gICHWa3/V49YqCS9mnCgiKZeFqTz0ae48Rf+jXNO2T52mEit+dp
KfQiHJaWtHoNHgCFUJRxkOJaMK0R+NOFr/HEv3SD9+Kv+YDNpurGsZLRRDnpy+uV
kXeo5tV9MV7CbAO+UKa9oQ0ACndgpx/w/m/I6E5aH56xmoqQFNv3A/HEM8Jo7vQu
sL5KMpD5/7HN6agqb9lR6BIKgElgGtA5Odk/3joRmn/MJZrgvk6Yvwq5cKuN5Nte
cN/yfcL39l+Le+2SSZlunDsJAG/g1ra0PwPLQ7uFlh2uL08VkaBLaQIeWJlY49Q7
lKqFLdiwHB02SA2xC5ys9EE92UKXP6P3TnSnQJufvKJ2xuVfYCNEwjB4VQEET+3B
hPaKVOnMBqEDLpr/8RTjffhtik2FLe/VlQf4kcdiZcHongvDNtLbcKvaqev31K1f
/zXUSfcEDmdr9w81UhWEtyHVdwmm57syPr8C61W2FDbXBilCB9e2xyT5fAC3Mwpf
RAPSK3Ds90kLVWGd42nVfLn3yR8vXk2ayf71rnrYodRWfsME9asiwBa0pw5abp5B
4Od5ZuGdxpqGYhwaJfrM0YoTnh+ErkmJ8Uy5qH0rmSQrct94LhKAnbIlYd1hKU1i
xd+8tQz+7+93MI5JjRcbkLH9r27K0RdL7N3Twhy8KryskzCSmxDnG9Hu1idMB5Tu
a1W/hl3eezuJIijDzpERAqj5kGDQekqhMwbwQ3ar7jOTUzcbrRJZAyQA5TfBFYvV
GAx/CPs4DllQYN+d3EKxFTNfFu7grz9O3gQ1ySoMXGZec8pL7oP/ijvTWOKVVqyM
6sH19XwICo1De9dlmR3OTVjXkeqAhLYWABlatvptCMyfUMh/UHfw+rfSrlkuQKwl
Ic+RRpoQxBP9PDKrKVwOq+UF3+mD+ncAxaCeZVztIsiA4zzp2mrRnqmrTmvrXKbB
Epz+Q2vpoBMnVAv1AF29Xup1JmOZ3uYsci3hLeoDOdmG9CNUT84kMDqHWS3DCdFj
8vA0HTJvmM76yO4IRpLfzBEFVf8lvlpcmAf75iE7U81+5SWUcTL0k5vNFFidhIYh
2hHZ+jOXVPi5P5ADZrV2Vb/I0ImpaRm0cOIvXGd42bNHIEbDtXf+0mnc89AjslOZ
Rz6KRWLjUzFvftfwKrkwuT6vTOBG7UtV9545tblsOWbCuwovUCnDF2+FFtrOIkWU
11xcyJuXlyhfdeTbqO21EeR2ay8XFSyelF+t8/oc/L+4Qi5UKUml3sp/g+15Q9m2
S+IoPnDmP2fYdmptZTH0Sb+bbCcewNyXfXOQVXIi4Ic+/76JBX5Yw8d5DfWUojAh
dqsN+6avgujHYYb/9F4HBc/sit8P8gZ4l3GU1AIn+u3WyBdhMPXEyNZP68BAxpxu
/QpTFh2R5F2zE7nrAq/AeV2l87Uu8uvmeDKxZqeSe4rPCsF1CmhT4RHb6a6TdsNv
Pn/H2IPpxFVr2c2MtUOpa+tkPe4idITBqkY2R+gq2orYhHvi4GUV5ge/0V3AEFaO
8lvATFw/AbsHinaviFenSR1zFiGkHNR7HwFzXy3kdRE9BpnYtkEh5eqkDzcYQgZ0
O7CSGq1cKOjCALOPKOZiCwXbnojRc6aJTxdXW4eWtKqcVIAkbNtSch7bgrWBu5u0
O9vGaHdyQcTW8C8yVQ2BaePz+Fypaoh5kpsZBPuIMSEiO8kqgJYHXdK+DtFZ5CFN
zlD1WSEWaAomVncESMLrE/zDLkQ97yD7V5+YSMlYpiX4i88dhaJCtNbMRWAv0a+I
Tjze1WpgOCnxAdIlNrFF8EuainylvXazsw2Y5y86SSNhWE5uzScABKgVvzAc1Qsp
gqvBjuSJu9usZVzeZD4g4OKRDJNdDfW9vaV1nTYzadkMAq6/PCdr7dWZlSXnralY
Bp8VePcxiDDXyakoYCk0nlxwCNE/ILwQXDWy8OvrZgy3+fTPKV8MKJFHnWAieyCe
aMr1tIDo8u8FHVJWOCJYqHNoCTPIps7iXOt1675o/uQvpxilIT7HPXnUn94J7s73
S/5JGUTQ3X2I/krso8gNhGh7dmstx/bU4AY7hixCVTi8YqABDFmajDJFhE1KaptD
6ggdBYY3qFxkTgdxzygooruLOpq5GVjaPlnBLChy4VYWFNYqA84GschQE1IHTmKr
dkUmxJsXShfNDO4afZ0s2t2pZZTJRAAV6+qF6/Gum6MLXlfI38L6cKuz+XXR2L5D
4VKn8/NjCCiBdoPqlH4KRzBUnJHz5SPrM3mS7Yj8YbF9UNlba6JYoRrjYxBA545a
Ub2ZIHYzbBAxoAzGlpC4ZH3TclNKxiaa3OJKjpQUD2ntV4Ixnrjr+axJ82m4poQ3
YM0JtvlUhPvyjPSZ5emFvohZItmj1TGh2J/l0p3wa9iMaLU3IA+81vaP8soSZACY
KSlfUdE7n2GSPLjl2h7Zc+3mXfF7f10q565i+G1qPA7Fo91rkYs2siACESLrSkQR
SnIuBZmuRP7UgdHGnrcqUSSeCZiVagtoskpbZQWRo+Lc489NBiwMN7sxpMeQdxex
CzlkVQ5Nk0t4YRLZXt2drSMnwKH0+cZJf2uQL+AR/dglFQ5LxTdx8XC/GSBwyJt/
agmJemA40wQAO6rfb4D4W83HrrePp6WI9Q4acQHu68kU8TsTic01bthJrQcWRQYC
wOkzpQ8nSj1Ys7rvqg9RO5/23FuExGKXXa1j5cYX2jB95eXHDhWtNY1uAowKMNH5
lw78FPSCV75KyDUSH/cmuSdWAk8PTfteROa1l+PNNQKGqo15JJEASU6dGGHiN7rj
Zm5bYAQCINogXltN8kkvj7ohtHpborvXqUvuzlcA7DW5Ps0b35uIPkc//l1ieMwG
6PaMrNxrK94zQbEGdCCOp1TP/sFrXIMj1w3B8ltnhr4Rue/r7YdIN+qD1Bf6cIbf
2FWnpRu89hp/Ru0ItmXTSZ6zaBTNn10tkH4nvBjQCDOWOblElTTaCchzgMa5aUHt
PsWDkeEWHckP4yIMzP+fn3AkzpK+ext0bdvaSZxNywOR+dPS1O1K8vOmtoRz2hvd
xc+OW/68w53lZ+MANUHh26kBwJ/JL4ZwSG2DZVtt1/iRoeUzFGEQZgkWCCyfWXXI
6Jh5lWMv+luOgRFLlyWIXRmCbmUEAU3ojwDnknQKEloFWl9r506z1yot2L9WQ3Pn
gFMxPsr/mRkNAXUmz+BcCHCdXWe793pLVRXF+kQ/l/uNV/7WRQurCEn/T5c4fPMl
zOlW8e4apJjxrBinUt8VYCcprSfkciRevTgVsaZve/m9yUDSHJmvEmtPKfmhsYt2
UrC0QielvJO+8vrxJZNIB5jUl6kobrj16g5SJNFIkcVnbAzFDLW/uaUezlOzces0
j98bWbHJjVWhsjzQ8/Oh7He/WwaISBlMb191FRrLx1f7UFyWWWukiqFJqx7sew4I
zDJascKzWq4oNyLwwauQyYgFPklxrBPwq4XoR9jmw40xrC26dfsF2/mdOYcrkgRC
mysMZn5d7sMGYZbBc5TSGoLRER1gXMdeRiM1duOhiwJVdVWiG6EzAszECfGCV2OA
XSYuTKC9n2TfEVXNSKBtILMe9MRz80tDPbf7dmPKhk4DwUaIomzvWebQ2SJXgZc9
0+S6jL80IMqfxEJO49jDLgvu7mI4pffduqGwEK+Vc00hZK5KtKhmUbz8HxJfy6V1
iE/r2cP8tqYSS6AWkcBO6tRI+9L8Ss++BFEfV0nIJmLsgG9sJjCrmdv+xKRqrQRO
YwdRvtkTE8Mw8leX4E95IsGsOY35daWfbovIFSKHOR6LTMtWRhU0CfWYFUO3DcLc
FLg2QmsrOdyZv+JV8Mj2ktXnV6uTWviXPmb0+2rR1GWj2COIJdlLIx1i6l6fcmEY
709qA7k7U3wqibxI8OeSV3xBNU8CINAgVNggNjlF8kcW9wGL6vDZsaMF2GMHsYgh
l5kSS6/KgCIe+B84U2VJ13b57Qumu9PlY5YIhHNLum57V/2L7UFMfSHwiCQ9ncZu
yWzARNEVjWU445T/K2/HNaZM0RWq6EOm+4l4E9wpfaG72PtUXE3iDrwzEufcpKg3
m2YEU6aFbpzRjkH9Fy+7sq0B9QE3iYm9FbHzgCUnCZI+Cu4IQkl7Q1PivT6GT1NK
vJANSbMIAw6B6wjH04AUV81yURq2Qsq8tgLhMZAjfTtwFtV1XhDc2rPMC2V9znJV
Qua9SdosdLuvLtiuPclU4BNXTPtsBuEiHaBhI3iIvVhBW/qnbZq8b/06yMfTUv8b
MJzu3/PO1rVmr30Nw2u3H3tayLT+6ibVSUJ1BWAOdre495NNrYp5NE9r617+LOhB
DaoZOwHQLvSol2ERIPe/gtsqJRzs+SyxGfneI1kdPHkQPkglfYfCivB+XGOytm2A
gd7Bg1fFCVUMwbNmx1JvMM+QAJOp4BJ8uNHkkrMg7pUN58ltMDAdq7ekjIHANfZ9
fqznUMmUKVCPr2Rk7e59rgWQp35FFHKEjq/aBCyTNOwWaQ11og3I4iPkCO/4KTUZ
iNDiEd57WH4tiyjwomXq3n2kc7ys2wuuahe7OQ08xd6oNU7mjnfOKPM/vjTlv6DA
kb1cQeF34Noksz0ZGueSSgGjwdQOy6Sg0NXeSw/9mlj5aQR2ahOSZUwCMy7cIMT9
eten1yJvoWgKfTuB+UQG1KXzZlWbsfJ29HhIiBvLkTuElzFoKAZFcecfqrwmMx7F
kcK4OsJZLJaLdaogXFbNcWxqYiXODxXk5lHWMo9CMP0l7Bp3VXQ8Kj/BWTjwC+Y5
wREBjHHxhtKt7JrYd/5GoGgCsUkMuqS9iY0kKV8i3XFBRw7ZSwvBqK2rZT1KFlTl
WlxmR3GiEEoeL50VvB+cm4V+aMfMbOoUo1vfzje2c72124UwlLjFb/lUjF/NoLOJ
ROo6nIYD8x8OAYtgs7Cde4VPiiQUlwCPqRNKEBWRTk/OjNaQquVDdDZ08idfFvLN
gBa3Tk4/ZNdBZnUoHTLCTR5xdl/7ErcKop1ubadAs5Ye9LDL31NjtOnygAsK7gcu
ykmpxZU6O6yjUYcjGfD/WjMgOha57Yfc/O680+xfMLZcOeEX8MQMSrzvkCX5K7DC
m/JTj5z6JfE+0tMrKlle3p0ugQAyeDJA+x5ULJtCiHqe5COpVG8v380vwjuupRK9
/dchDrz1RJs98zszKgKN7ATf2Z5524XOnnG3jbKKe3vZZU3f/v438ejd3JWiMjXP
pzhGxT/i9rgwz/duhamzOHKE2KeNx6KffkRaXCIhv7Ojm3EM1jwL3CEqmzkqbH0Y
ELzCGF3hj5serwSmWhmkiNkDEysa86eH6fdwQOK1AhWUy76JkaYB8rY9l2yamsU6
AFSkhpHqDyR9hJsgrkAteW3KuXW7JDA814fUwEZCLhSDEKqvzX5RITBXdQ15BMW2
i7GegtOclQLA56QMM5WYeREQO8DMcVW/iqvRSFNgJDypCBOHjYI9uo5QpLrVZ+Z5
F7hioTGMY736ndK6F5dNtOIQoY363gSdm98Gis3DI2StUspEzpH77V8XgEyp5hEL
d5xzWJywtpciI8oqynOyD0lXEnlR6FWzQqNGf448dF+mg+hgxcuOiPbl0/bcLIQo
QOUm9num7bRG5W844qPxSVNmcecN1KCEzfVC+aTg6XIJIDQZCyaYR/ZLQ2XquJHD
cXT+EBgALksE13OsUrfKOvxBOXyaeZ2cMPDorwxP9QKn6vMhvt4ZdtkQRN/VrgxW
sOw9oR1cbl4foBTGEbKRb8k1wJn5ATrhS67FAnI7piuUbu+tRI6zDgyYvm10K/6Y
e5vUMJAMlCktOOuTwAmSdg8WrauhAehojb7+ZfdAnze8Mk6wbx+cZvp1hqlGSpnq
G3zo85aZTKfN2YthTMWzHqqQer/ZMWvD3B+iiADA+OFhuwhyDpmiEa8WQI7HcD4S
dOiYYVQkOYZM+cMVGaZg80TmZZSHPkdL/dnVZRg3xUnAXcec0WM+SSqLqS6u3ddm
Zl859i/ffftKT8VUO977c2m/PTmoxxpMby8fs0GMdSwMMIXonl70MI7Nu4u6ft9X
nGl5jgUxliK3uhqfKDp7g33Vg/5HSgY7GNuuBoBAUYWU+NDLoYGlkKX9ndmu/fYH
HevY7EgfmPaCBJ3Z7QmSmziyU8V3OZ9hQLJn8VVcFL4tWozV4kvFzESV53+6J2Zq
9PVoo8TjeKqFrQvvfo0H7LPTsGcXfY1XyLvX/Xo0ciDAS9tDih4D6nb35so+XjMh
mluh5Rlt99bQwHf0A3+jkNLRaMWnpwnDsHw/9mJKhwAQHY7Tn/0ixmwNW7xRdhuh
GIylLuiM4u/n9qjODBcWc3U3t5EBNDltIo3jY7ZpVopAJqU8056myCtGjiaGg13d
IHu7x3izYjKDkx+xQuZLj5hoJIuaeY4ltDXtzHiFECNkhaUkLiHvSSTTU3wMO/kJ
GmBWUavUiKdQJUKsvJG0y/Vp1rYTlQfJcGMnoUIgTIEc52K44aFvWUratjj9WrRr
Pa5sieJwDGHb8sgLCxydwOT5d18yVjkc46c6bau0wG4h3ORIYt57jRNp9lSAmIoS
KhhCvyy3AZfod0E5LLUGyBQ73JML5jnRLgVjnRb8jV2CRBbP3BECjuyRhV5CtV6N
f83Q5UfvNe/hVYqXhWAkeSYcO96deQVm41kwmefjWN1Gik2DKl4eAn5p3ok1pdVX
xmb0KbC/K2zaebjcJjqsLCKrtu3E7NzK5QPMvpFrWyDL4A788hTvBdiyqE9YHK0c
0ztLVQ/ePE+h/gWa3/6LWWz4IPJol16FwpbcZr7XMpdo/55lJiXECLd4OBcAJ+tY
1FhSSULGpmxKMtZ0KNxpjDFekBd7hCt2i53lTgm4zDto/bPkE5Xbx+NjgdOj2Npl
eYTn8LKi4hvhhswVCuxHCdAD3vYdM1I3k4Fd6q2xRZrCGIy5tXpgYuGUiFpt3Pt2
oiQZdRIAnSf9BA4m5KklQPQADJnTysnPzH2j5gA5c6IuTqjPoUmGfloy1OXVHRgv
YYdBpcpJf2GN7Tgi3EtGqSq55EjQyg9A9dqh5ARHON/wJZluF30icZFjVwPHOu9w
wJMXOQkjrTMUQ+4UVVbiaOVhI5qdJ9TsNLIFF5K6/KJ8AEnDO6eFhpGKjvIR14r3
DPtojvA2S6H9jnLPx8Nn8TMsWyBjsF7hCqOeCiMEnTKuUJg7D4zexk+UIWjcNeyE
gmMTbooTDSc0IZA0gdmKgkv9jwCNjdnDp3kdmasAKdX44vmLlOw5ylyW2yi1/9IG
ObgprCKYMUPnuAqgL6h0l4taaf6iMfkCc5suIVNkiDJFdlkakuy74HgxURIvnMwg
bM/mhoKCLCGKFLHVI1VycRH4LGwyd8P60kjRcv19LXfN6erbXVd6F1mNcFPq+QVg
jGPjwAoLGll2j6KwTL1uJ5pKEjxfF3cTaRac9/CrsfiiHEmw6RodnHNBWs1SSKG2
FfutIPe5ZuglC6bEceTWwM9R9Z8l6WsVBAd8PE6X6gYRKpawPZH6ZEfBTvkIP01a
uTn19nmxyZxJ7cX+uYjWyYcQZltTELfttTSyCkoDVK+6VyE7gM4R8Anf1kZyIzm9
bt5n9pETlXXqFkVgdA4gABjKf5vvovWFSYegICCtydyrKmnAHY5e3HOiSzhuf+eT
NEtW1Vn/UfmSRuzJY1QvyNf2hbvAcO05BULipeZmqsuNBi90800EUZkNuPeA77xK
DFed98IZI8wW/MGqaFSb7olpjjC5dpKc49TcCTWhBH6U6ZLjCn5wIWJdbJqhZ5Ks
RhFpTxn97EH2r+iJqW5PSziWtx2Xi/a16zUW4d5aFzX8wF/nDgC/yufC4bTvKaOh
PFJ8dXajBH5lBsKwh+Lc6tQChCBM585n0A0OTF9lY1ySfz9Md0qGZi24GkmG4Roo
we369vL+zrNyFav9S6zVwxuQluPGtY/UJ0BiIJExQQgVve5CY6KwANOeGKI5gfbh
Zn8/G5nnV/DL7y8cR89j4Wc++u2+90h7QgUvJ/ksHccesM6wRZ7PMs8m6zzLON4G
kKEJaNfj3gJkO5o49nlebKAX7mhhaqnHFRwl5fyrcy10oEw/zH9Ld7BuXxkcy/YY
36C//ANwFAnVsrRy+uhHFXXYpkYv3Hqvz0LCyarYZ9hVvQez6gf75Pm8OpJaMnpk
85it3gqzkswfuyyBhjQhnBvtfett+DKpd7hL1ZBkJlGWQRMfQCBF/luXzbDtxanw
aKBq2uoWyz9a7aC+1+uByeq05MkS+jWsZM9vSJi7bXVDQyndvyqkhQKzSMKneM+4
I2prgoeYV1hIVXIe5YD8DTDGcjYwAvoJ0GNnrnkfcafqlARNFwETPdGwr+DBOlyE
Dyc9iYJK2iDStB2g0SNs56Eb4Zx8rgNYDgHK3oDOiiqhMjDOTKlue4VSWjz8mCr6
3FGmATVSu0di8p3w+hjh4RMwM5BrvMuQDry7N5i0IYMR3O+1RKI4ORDzABUD0t8d
ORiswd531SjZUgI10VlEtuPJB9bym2dEv+xrBQLSiKfPfk3bTN7UZjahjo5qhpoZ
Hx3erGAGkEOjBZ9/VitdXbNVRbAI87uCc/GelHD5X4jUEpGu2ZGelcEXKZe7pbvL
eriCUSSBpzVX9AMQ3pUi2CqkJhOe21VX5AmteavgGd0GKINiSEzPVYz6i4twergz
21geZCH776YNtxaIQjOXu6Aoks+syksgm6OEj9Qff7V4mFSbgX94/LPFyDrCPtPf
9xVNUOC0zC50wJlP+N72oDc91MVih+eZ6iphUMXYrdoJWkGAkSy5sD7Ai9j8SVgT
4Mrnk/5wAE3rhYaftB+kx6tocY4e5hBozjMSB8dHfh1GOrZ8VjcSSJK/Sl6fHyM5
DPFcybqpsiIFaFacX++DX8Xeae9GOZI0c22MnDvq8AamkfS5PuxxR41SmsidWMg1
5eDleJlql1THZNyBYTbvgI52jtDbQV+w9sQG1rlIDO4KXG+r2nCYPiOHVkPv1D/S
EmaZqT9mBnAPbJd5S0mSSDiwjieAS0MH1hkSGinAeSeK6IWB71zNc+z0+NODYT2L
hEF0GcWF+7tJfW8TuWNw40kuvJZfyEVMKMjYkLi9S1JEoBy9nwgYa/GmEG4IoPzR
A17Oimj0dWm0Rgh1IYl4i/hyfnGtfXHqOaKitwTdNFVGCQ2E7KmEGNCRuu0YQDAh
9u+QRhj9dF2Jg1pgDNEzq1xXnx3gwjfg5Oy6vnruP+OsriKrNY3vjTdGDx/lXabd
8cWOvG1PzevgjVm7fOXe60mnh7+FnSwmofisuhVrPqpbw7EWeJLcfVZYH5PuqA41
XnApM1NdDYpuX0AyvJFpNZBO7Psi3LFZZRNPT5eXdzS+mYaP+gb/BSweI4HXn63I
+IUxx+3Po5hDsdMy9BkMyBpr4jD10WV4Fvfg5dgO60laMwwfQ5wzCRnX2uTm8LQz
uWWNjXVvGd0RML8qE5T479ZbH25va06PxbkUMvekhDpa9dH7NEv3UsV/px7ra3In
4C23c6qkBVy/59EjyupPT10Q5DL+P5WKfWBIYaKS1QiTqO016/Nbwy7GLzFKHTQU
ey6aqTmP7464T4Gh9YlOGs7jCjIQ5MhWaodtYC0nPsYgCU8nv/HoSi1EGNEu9MD1
h8yTZNrDtbwHQSgbTYLwc+SrsMp0QpuXQL4NBeY5XWoEu5/OHYtvesr55+twH1Js
/FiDzKRar2HTXuhuVVL8oEFwdAfgMAEPkYcprf4kgtT9arvRNztyxHbpnH4YGomy
8yVyrOv4aO43i4pbL3JwbpqSFF0mtU5gcSsYuqGk4hflF2fXPfXS7q3H0TQZdP5w
PJw1St5utk9KeL2EollqLCqMvPKDqd9pSTf0FES7OLoRIUvXrO5dwEDzCBCOWsv3
NFWHwKvguc5yGoX5s59p97PPam26IqdHKmux9u0O9ieVQtiO/vaXjcMJ0OMkzuuX
RV3iNUy3C77sWcUw6c4wzGw5HHMRWOmZLDwsB6jllfleivYiuNL7ArLP0jd9ieJj
3B/VZUHn0KMMRcYG6JaZ9NSmZJS8mxUUQM0BF7XiJx4smDM1vhQIk0EX7Ivck0zr
Kd2yU3S7VRaHY4GWqQA34On5uuJ0AwjeqYH6KDwhwaqjZPXch08QDtvsXTrJjl4E
EfSKr5Pj1Q9YOqtZB3lucxwZHO5giTzm/jc1vX5HuNkrsgVVY4rLp+qnLqv58ST8
DxsZeVKHSMcbA2DINfWODAY4s6peS10e43XMH1todFsIBchEMr9UqK9pR//Me27v
CNtd7g3dGDnDIVxFeNwp75UznLm8sMo+WvnQfKkjK8lgyPLe7rdQBkWM/6PJN8KK
JqSEI38FDYY9xn2oa0S7bAUWK05UX+2qAIRkKawyQ5S1mfEH1DO1syJel1FH4fuw
radbkx9u9jQirORxLOgq3NKrUpdV/lZV0nHSmjDupEaeQYyIfXbXi8c6g2e6TXqD
h3HlPdKf6j+k4GYeJvLHQ5DdlO5R35CNtI7O+/zgsts3J/lUS+9t/n3UNS38AKHu
iDUOmruXHzPcyYQe1KlN73NuHhnrRKjfAvwnGryvlHbaTYLd1hxZOe1hKpwhy00i
eaC1L7NgJhl+1YoZbpN0WCUURGpNmmibF0/FN/7WWIKkuObpsRBte7sBQQYG6z1B
aO/QjIqaAaZr/oM8PejCQEsIiWy73JPHu69JCJwzc652WcgMnzLoXn1QmGcXHZDv
wcVddeiiE6TWI7eX3Gezkxz+bkR8DS2HVg7pc1y8x2S8tufHiyV5V5UBaCcGOWgD
7ZhcGfHmFmVUwXaVENcVFZBIkA7S8vK/EIlWXapiS8uoIGX7MykzYYkgabuKwxBx
cIAmbCWo+cZ7+YPrTrVgn3miGzC3hu/6Pa2drh4eQfPFz2IynRV34VKEbdfUwHBO
hRbHIh7AJ1Y35jjbQIqn++cNVkuQNH6W6Q7eIFPT5IYrgazjSRlEdwL5o5HPMTdm
pYlmOb2xdxFAOP0HUUaV/bebfhJkNIMMO4CjPN7SHEJ5IxjK0Nb6r1afMAHkQCk4
iR/OyclQrxUTK8X03eTWZ5O444LHp9Q4aW8vSiLW0ylrpH/sp2wojr9K5JrRJpL/
LBx3MAkfZzH5hfWAn1mTujwQFVOART+AtRXd9DTX0zz7v7AhuGSardc7QCI/0uWg
HKg6+Yyp3sHPYhBKw5YnG3wl3N8e7j37K1DjnRm7bTjCdxQQgElvVupIqgMoOM2Z
r4DkCemxSjPjD8Z6gCfR9zolWVvfBQXGpECKNexgPuMJ8Ycn//39GvCXukowdwPy
8hsDVYuzTs6sTqejgYl8TIhWp4nZO3pzW58UECLc4TkODGLXfKNjubHKCOxLsitL
ncGLVd3l6subChWj+xT87b1J5oGSIfJCD68N3Ju0BKgAdbwBie01+SxNwQ0QIFoC
xzfgncgTCBvMKHJp1YQAKLlLQmXCB0Zg8mIDkWZId+BrYlhMKCQZzvwUjhVKJYhH
ehfvYuy0n3oD3uH6D3spk3H8xR5WPL6+6Om05Qp1URDTb1tGeboraoY6F4sxWtRf
VMM1zSM4EZRpaUs3au4hvFAoWZyRQoQW3jH5e+8Q2ZsjbMyz5AaKQLnGdOO9tj7w
NBmt3TPIziBx5YgK/03GXf7jXRzjcQ+zpTkMw4lcqFSPulNXEpBjDZNLJuoDLWWz
uv9iC3ggaH375iCAo+0WatOHuTFxcZ+3/0Z2lm9M2epmIIkgkpfKuRGIGjql4xG+
R/0Y4W1F6+nb0w++odTw4ijHEXsRgxU/JRAJtF4e5m8LW2Jkm9cD4YVhzHEWyCUp
NevXbn5VYUevjVdiY2jiE9PvdAjBbJlLep3wc4OKdfBg6H6XskkhhhhW32VjhH2T
eSeGpvWylLKKKKtm7vERA1Q4DKwp2PrxcVNMZpol/I3XfIL7vOsT6Q1GYmXikSVR
ROreQ/B3Mpyp5enGRHTVxBlGfUu5/pyGk51kkI7h9wpqToEWszkvnGO2yhla+JaB
QsQhpaw8S/++d6jD6moEMz+5+G6lRQv/tBoJ089YtyNbyqAPDUB05t+Ndv+vL041
Bml2gFhuZt4+X89RBzptVMKAiw4HyygRAisIYiGVGKiswxoTtuHn4mc+ohLBNG39
1MBQJ00aNCUMgfWEMkwFv/OcNsGhFi3XQNVyu1wJE0VW0U9FM6Mesaw/g0vTvyeQ
mC07xK/LBGwWIUpA82ZBoP5tmJn+2IxCirshpHazyRayWKNO8SR4Ehd5qA4sEP4s
dMKbohs1Teh58JH+V8lCd2bCETFD6FegsNoElGnCEMN4c5dsvQLfGE4R8KxX3wid
jQQY2IqgA0jopkHAploqunwtMcTGp6LiLQSP9rhUOZF9ks3pbUGd55u2APVKxJr7
T8dU9DNKVs1tOCdtaQgu4Ryace0F6nnGeF7ZAia6VNhftrxymF9ChLl2SdrPNNVT
W7OfYklTWO+omH7Btqfw6ysJOGc0p+e5wLUSc1Bf8jpWsRrG6pmFplvUOsPP5QRL
Lf8Vxm3XAY5E5y+wBy19xQNhO6l3LBgNR23T0nI8ZMFIZ3Vh3+fM43hwsUWHaw14
XUGtyT22PXRcCxArKwZxxjRn09yvSmWJfl9H3FVUx38riGPTpDQu8o6kDFwy5N3x
CVLX7YtndtWYlJ16j+djlNu9tL+4dswlSgp69Xm/s5jacvmg5nIoCcnHSrdzZPWm
fo+VL221kAO9ybSbCAKygRQEd5wEpGfwCYLWU8Aw4I4k14NvgdbLrm3mBKqyenoI
YGjtjDbEz1uMDdKIyaL95lGXUm21/VNa+G1nYbNT72+p+hIxtHVGwBxdnyetzL8A
B8JNlh2gudfnVCVn30xAQgMsUsmrAS5fI7IRj28poDn9Ey+KZhtqImEH8shendfH
SRHZAC5ViOZs3LNfZ0Lv/QNQoJXLDoIrt2vpSfOKo1yzfr+GIcK+LvIV0bfm8wB7
DoxIm4kColGBEn8PIe+3tYBR4HpQbaBYuk6k9CyXzKkLaGy0tnBBGlxRFpATG3rZ
pZ8B1s7PsUPzjSK2eHQ2Nbqg9i90qSDVoBRF8fUBRm5s+nmMxTlsO3tCnNpkl/HN
CAB/IQho0g/Vj89dDhqXi7I60aKdcji23A/NPs2MT3HIi0vSTTQVn9YOOBnF3/eq
tyVXwGob6iBsykLZGmWWCwQlHri1s1XmkfgF3iiDTX5v4IoHu4vFkZwHI4lChsuS
iXEGo8ZkmgwRajbwIyp+T/uvtca8nNxWncMgbfyd6ORZwEaT1OvFG+/8k2jpGDu2
7P942pBubzX2HjBkuSmz09Za1Me4dsrdlRV8nFqqDQjw3zhrU/mcMu1dPQnuu0RG
2S/hG8IMc2/3aDwQtAzQVOuwVcTIEkx8dIirH4L6+Qy+9uOCl5KIzwl+B6G58XcO
xkByaM3QJv7r4Kx7twW19hXX0r7onR/KQpMFy3hlEABLiClCCDcFFkP2wUbF9SYP
nCDarru9i4pv1exXPtc9ny37iH12P4TzICt+78dTOqlKbjUa6/3mHpIVky5fV/K+
8OitmqDMr3S0ItB8+KSpIjIdjUbb3kQMvv1nEfXhr8B6Nwflyeh6AG8FACrd7WPv
BP8FCVme9kF9tvZh60B0eX3VVY48qTpzq0hr5nRcQL2RHuocXwFclX8pSoJU/RkD
Dt2zYpBZtR8X/0cN5Swyg0OdI092NdDpAcJZpA4K5+yPkuSbz1rT59fpB5trkMyE
DTqyZyxoBu/z0A60W6susGHLhAHG9fVqbAgLXJbsQZeZrIPb+gpWkFXwG8R9PQzb
wE1YGmb+XobAl2AjRS7v6Kb7jqcsVTRPHcmQ9Be92lJsF8MT/28GMBko5qM6k7tB
aOo0RQInve07VVS2BYG1Imz7H4foTnr//sktyPpLiTvNarE5XNb9KN7+VNR1LgVl
a/33VUDS3bttYTohsfQaARPcRKDr/Ayaa1B/YUFL80sKdxf/9m9adxNyPdjm0NF1
2CAQBLPEUxAX86RNccX1lfskdYr9jhVjFCsA4tRqfgXwBps8bkf0MLvG0JJIHp1r
rXg6G0XyP50/011QauTgDXX55hQ68PLONlesA9mUjloXCjyj6BTebYRxcGuE33qL
kXEVJFdQ5HFP1cxGop3vZfIOCXG25piw79eWpkkKa0gKlntyfjY636EjrnikGks9
6kzm5+wkMDoS8hT5ogP7shUJjP8JBpt4PJPaNIL7URZ7g+ejD/VkFUWrFfChzV0F
Y7TRS9xiZQhW5rv+ZgHYCPJoPXQBF3Pdd6srsxbuH1YCFO53aLdFZUkVTUH3r8pt
8EBxqigKIXME+pkZv4ol3b5iB9rYjX95xtRsA6FLvShUN6N/dT2ZLA/Qc0E/mBLj
3p30XvUP5Zpwfqc98xT2/DuKT9p4BvmBX8hEcH2xCkGdyC/t7tiSKqKxAAuF3tGK
HRwddAhGKJInX9lR3+rbmcw6QRnkIgteA7XHjMi4rWCl4uj31YeCVnOywivLgpw0
EXRrlLUOMYuAeIA9hWiGmk6x7GcqQB+zhqt1Ag6Ddsl2ZUUnSV3n6ZBusz0v4Mdx
BrETh9r23kj4G7dCoGOmZkCASlZDnZvpOVvcSV1XdLYWmF+CwFZAMN+L1RvZAGKr
5FSKmgWrUQfOjSpUi/SrS2kxecxgIeAMnDUwpHfty+hOHTrTKKaXxm+bGMgwtVKG
M7nRl2ecQ9DAqwTCePXISPplOXWZNTSWO+qzkrFIAh6Iv+nxjTO2fpi5D3UxXeCq
cimwoAqHXO1O0nz/l0Vnyxjm2HOPv2GtlJHTocE7SNE93EjqUBDAIzgQsTrj4DeW
oiSyrmtOQAKxWMf3uagAfa3QeVZ6NHG/HL+hu8rNGOAlfPj4V0UKMd0SqM5drOCz
BScHX7Gpxi3d2h/TifNCfw5B43awEDA/pMS+1ebJYgLHQE8vs4Q0I+tSZt4wCUz+
bnEcmlEDTsPaktvIaE8DIaPDf6PosQ/CMobIirOoQiM/qFVFzhvk68jd7+6S+hwD
Gk3UkgWjaU69K7UeIcQ6i84M7RoADUdCvImbaWIcKn87C1FJwDHjE91JO9jahUqX
k68oOY0HvF8LHjMiceRA51WnCxUrloDmlawaFGvWHpcwIbuW3DQsBMcq63vlLJvL
bc1MG2XgwEkl72xi2f9iy6MIPNrbvJf7fplpSXli45RLiLkhknlCteJ7yZOJiX2S
WGx7g/Jgh8+TcoENRhCIGeKpDpgmi72mMQ7cHfPpDN0YOl0yt3+V0Qemigy+7fwl
kURCgeo4WQ5cw610HxgyBtKxOvjIc7wL89h2n/GU/UyRwZpkh0NX1LPCNLLusTUX
sor5gdrx64wnysfeiCmnh6UF07J6xuUhVgz7/IBGfTyuhoCve9eattpXjVhlStS+
6aYT6RjVUBGmYOHG/eOGk6Q/VEzp4Xtu5JCt0t7NX5yecxGPb17CKBLKqnGQgrup
r6BtFXukNLOfl5GgUqHUUF11emztK+JmAFGbwDR/N77Fdge+44jv5iO/60rj1UZ/
NRbs50cqWRo/uG1SPthhAiix6DYc+gWai+iauY1ujFr4JC+y0Lka8OgKPFKNgsSn
k1FQ9Ekr/9v1ML5dVqrEBNwAvkgyY4ngREMw2Ax++cr+OxbsLpMj3fXnt7980gES
gnU/9RP0KC/XH7gorlzxw881n55F9ioabRpFyRuSRX5L7RNJ/zXn/EXEkRpwiV/I
beNbCkZ6zYb6a3kGaru+ukHk3l55ArMTUKmpwoviOE/RbD/RRA4lUGuHAwjOloFq
u+qW1mzCm1aze1p+2bx3fbbxA5ld1OSX91HbmWvga3IZuS0BO/uzmXvJPZdT+leb
va8fsMvNbsTSTcPjN4BFYyfPYDB+I6aQRCMPuyTeTInVgG2FS+xvdqzCBHy9LKPj
NsOGenYkUyeI4FAUqNhYeEM0Nt0KiSl+JaXHRHlyQkDjkJ5F0KGoZJAyG4WIDm+b
wY1zyKS9WShygIGQ0RzLC9jKkAs+VcVJeZB6YDDyKX+pbZeI4L9FkmsCkp93CVUx
0AzvTAJxF3U4mVYykVCn9yHvkznRDWeCaqV+GKfN9NiVm128B1nOlq6OtAJdG20n
NY8dT7B9mOWbK45nYoS4iBfORM3uSNgbTye97vdDzAbJwZ8LzR2Rf18LGGO911Pl
0abNTT9ym9DEGjVi7/S4FimRsHq7Me5Mg9II+L2GifAnaQw3iTJP/p2MkLa1s9tw
dKPlvdRSRXVZM6Na5Ab3UsaJuiM8xC2gSF0qKijxdDJLDMY38f9ADhiftn0JAaQk
KnYLc6XMQ1Pep7RQIt2aTgOaNnYEVSgp5/JJxA2eURpg0REMv3/yy1lz0L0uWiiS
XZ+uNtU9T0xyudYxH46c0SmSYVd13KXGP7oph3+Cc9cj/ax4iRRMHWcWq2HiC4+m
0KdcexNfE/aRKQG/N1gK0TTegHi0cLgLXjiULPp4pi5oXrVRjJucTYV6sr7+fH2A
v5vjCefqsQxf96K8XBlgMmG6cLHKstlWP2ZgGEyOSKqusaOurFj689GJGZS3SG6c
FuuNm4SP+OW+jHKazxqNstXHTF5zhgudSYEZkzQm6Pd4EEGmpvzQ1uVHc/h1U83z
op3VG1w8VaHe/+T/I9+3cS3LqYqgc9Z8pGrlYm5erK/eSFpf7naOyRDBCoBOV8Ug
tTMOtl293XPDn9IWNeaOl0Ah1OM48QlgTDMA+d2PN7I2Tuz3cOiuuPcYNbOJhVJt
TpkK1u7E0DliRh+FiG6glKKCvnnhvsb4Vrh1eZ3sCDXY1vg9aapJQ7PIVQxNpLbm
vvl7d05QVFDZK9Tc4SIcmEpXIABVpiqkxLg/X2remfrmO0gauhQviMTDtvPRRNPo
gLEMTZ9YAp5Tj43k2P5yp6jKZGPkN3dl+pmbtk+mnHIgPg9+QwkXOiXut86N/bro
zDoSTEntJBqQ+gaD6oiBPEErtitJueUg5nxcQSBEYiH97ySXjy3jxHAAEmMv0D1v
4PeclpZXD3Xkae58PrUeArI1paRoU6hrYqyLWOM0hXXDmEI1Nm16T0g3qvcKO7sX
K2iLtNWJxoAb5KOcLA2p2X8prkCIXBdJjFRGQG7zUrrZ4sCo48YD6fO4HQWwyRhc
Nh0CJjlP++xJcXmI/M1LF3czc4XUOfz9jl8I2p3ZIqNIkesqADiJwI/3ybVK1VL4
XCx7jr/P+N2UnwAf/263EVw+FsH5sNMV17vR6xV2yNqQJytPKlDVxCcRe6Kgk1xB
2Sl4+eqnaDMpGcYUHiUX+27Ttx6NRhLFLwKnBhNkrgZbjvulomOOW/CwcKi/1usr
c1J8bPesbzEU7La93NTUaiYtu6KnzX9FV0PxK6VwLWMGsU8Y4hK0c1wL0VQIQC/T
uU3o241WXWswaYuLJqtZkmUg+xV1HmgvgVPzKVARC39sqV/mbDKMbNcUqaXAfkeN
0KPHYQHoP4U1zPnrUwcDmc7GzVnli0Q0WbHrSVEIwVuy2NX/P/GC0J829+diJY2n
qpyDh1vgRLtR/AGkNxVjUErgNF0duvPwVNLvE2cM1uDzx6Xc1iEO9QgPu/v0kptQ
5F5bO1J5K48oh9ymCVYxadVdPdNw/rsGUPeh1xdTotrPVt7UQB7eLtEC/SJjIynI
2q52uPKpTR32Okxyxilo3/D4uAodBdJRE2MQwqg1u3CzvulGOmV0RO3sL7UsaShr
O+xf3K5ziDu7d3+0YXwlsefhDxBHNnHYhKYKwCLPYsNTqSgTZhzfdgR+Dc52ZGAX
byLeKtA+i4L7g+2XyIBC6yf+Sy6J0FpUMrwkuVRX4LZYvfgNt8qlxJHrtP1ne2rQ
DFQkInoSGScx2Yj7pX4J3x6927qwxFHm8qum/pY1dEdrXGVse39MDHu6QDBtyoIl
clGspDf6iSPrueRFAXEpFQj2hvcxwgxBKjCOfuitNRRvFN05UG5z2OrTQPZM2XLg
7NnLXxWcWFXMC0iC4nsRgys4m9FwQd9CkCH6iT5RJM1qM9m3XCZU6j8+EEDCV4+G
YunFfuZYTKoVCQhI+GwSqhIH9K1Ah8BzzgeoCQb0//jEOOWGLXkqwuv8NJlOBH4j
CjdkQPE7PSdsZA28TOW8QZZZQ4zTEgi6+2lUhXOVSEOiXrqgPMRcjoNggfgZHHhq
I80Q+oJxJIjRL2vGaSJMwc+T3YqAypa/9lypeVncJeojGrqTsPa4fpcAxzO5pD1L
dCkX3S1Auj24GoY40fu8U2xOW6UlcjTuURVYJVX3Pfo6M8uYQEhF8WwO+f4uidpK
KoRXswry+C4V67jTlVaKALvMxfjFN5RRm8nOget1F84FpGrewDuXcUud/qXclKyr
hvAXEK9kV8AvyTgmZhLuKNCVvkweLpAMDqkMpweCnneNsRfI1s9hz60MxVSbz022
UQAONaKnG1W2J4hTDZgEStFx3SoNcKUyfzjuBG3l4JekHizKe2e4IRa5zX7ECu0o
Tr+MHIBdfmXgR2ykpsvYe4aySAwL1xywq5VsOv8R3wV1MtP3HBD18m1U8NwY5HoV
GYnqZV+36jbWrWE2kdf2hnsOKD+BVLR4KHK9miLGwI/iKQj//Y72F/T8dJmUtnVn
OhTleJwXpkJQA/R3X4aPRrzBrFADETDHN+wXSNxPq5U/ClfZ+omj5kVcqnUopzN4
dSaSEiwo8G4h32sZj1D4Zyaa7K4lcxA0HRkELFiVrhe056jz7cXGJ+gR7VvPPiKr
sNPw+U8BToJilIKiFMR688WVQdre2/R+MsCNVrrDsMfo/3ypRyi5/JPWeoiKhXxz
t054nZeNRXBMNIosYWfpZiJCzs/Ha9tSy5jHlHhdToa0h8OJl1RJiqeDHo0WbzZf
R/6pTbQAMzx8IflU+DztOp9Dwqw3IMbF7niXzJQ48fgXVexc10CK2aqlx9I/NW5R
2uK/AucckQscMr8bt/3kUQmu3bVhp15/nq3pc1VQoiXTNqZSSlZ5tP8vPVnHHW59
xC2YReLVzT6kQXppEIjvgCGmvan3buoGcVBTyljOUPVL8UeVgOxXqhQ87eW4Dpa2
cVlPdhLJ3gLfp42BhJRl95G4Yp8h3h82RZCbJJOOYq2MKogo8dFb8bs1BkDCVDE8
xE6W9F+L+UgsAJrHPbmKMTecW7Jie/SVsb93l8SznE63vy8lXn1rOSaU4gvn/nsy
MRJOGL0RhxoB9BY96INHdHK++bRB/1LcqD0eGzEtSFbTzAkwjdvL6oZR9hQWNKxf
Y0ypnGeqk0PkI4ysOG96Fpuv8Sw36M9/TaQ++7Fl2TZYJDal/bTDq3B8M3ZhU/mS
RkvXAxOXb+p0s534LwzzHt/pihHoz/azh0vn2+hTuUtetnL9HZt9V1hLKj33cLa1
Z3awg5tEPdmbnxe4YhTtO5vsc9PEx+cED25ngkiLXkY90TK3rUZaxJ8TDsDkOWTd
eLaFI41WrKwj/IusZ9oyXO/gbWrnr6bdenvFzuSxitfd5fvZmAe7hL2IQ5qgdVx8
Br8+i/ybKS3OjTzoXNMDvezDJngoHhUWhxKCLJYkd+ItFQ8279uOY655KJc7zQHh
/g4+GnJaMvNZVBOExMnYhS6xenpWbZoXJLrHB4J5KgiqW3f6ZDQ+mL3jDs5jBfPT
OEjGtVc8TFpYeXjkslvSO7Is62Gc6aW6sN9WVkrkbXNnyIXwLtJaJw0Lr0sxN9rZ
xZTCuGp7eZe7tIlKz/JwLwXBxkbM5Y7/+9Rrd825+7RlDGlW64SwPclybI6zI1vV
9GgGHYU/TV62AX4+FEWjzMDOVDTtZ7h+xGS6DkKKmrM147H0I1F5ZUwog6JjGSEv
EseY6SNJwkOe5bSwhDqKg7PSQApMKROTnSyRRn4vCcC/PSnRQCdgcpUupNXQGj+b
hPtwTPy8pR4UOHAfqJ0dcSsJOhhk9pYe48zF5D9pct3Q3w3xuiAmQDptMUG6CL0m
SERv8YN45+vhRv7BSRurpg7ahgZqIV79JcRVa687solzCxqtfM8xKwoIEi+OZXMd
+SYIDwZb0mHm5dL1Bp6HUiu2Wq2Kpz7XrFmN+GrsF39g+UI/BlyVC7EKW76NFyYW
PB5YHgqv+OKBrrNM9CeA9Fbib4xGU/+6YnewfqqAWrzZkuWSnjV+66SjX39bQ/3J
GurnuiKzkkTU1YCi7WeBHbKgMXPVSqM2gWWp0W39rCKvV9TAKJ3sT0Ag/p5/nbO+
FPlvxVdyaPNfG5sDAQfqBaPnwO4bpM4trtrayKraf/JD93tzufaVWPOSxNDVJxsb
e+izNUtoCX2PFVrdYpvfUM0M7PlsTMRT3MJkaWyzDezFmdP9JxH7z/vS4O3OiXCf
OpnE0nByyl8M0AakLesjSLkj+hg+g1Wj5Mjgx6o1InNOUPAJrfIoRCHWM8WfdSH8
+VgttDnRCiC/d3qa0hTl8EKxuFDUBlByP1Q+SsPUr3HMv3zth0+t6MMdPbIImvfp
Tpev9fSGTEY5xHUNftjqK4HIs5CpWRlXg28Nha2nVA56YlkkkRfQ6qrSvTx6zWWl
ntyNvQAhXn/qGwGQw/2fCU8hYUifl39Se/P1e7yvdz5MHBWVzpih6MZpnwzfdefq
kDW0wlHAo1FYdgZWaMb4s+GcKcCIF169TqdplGgGYkj58Yci3HtwqyWjNwGikVQV
Llyq/0jvl56uLOQynrE1vEVExSY4tkcFSYDFvifeZFNsLpbMYBxBQ/O/tS3eiG2+
1iN+dPle2iqVDkAry0qSd+hsHl+Ue7uZIPT1Y/UDv24JhlC6IXulCtCBu9uqqOPp
pSA4dpbxM21hHwkHMPgs06QH0jE0v6iOrzafKehewkocdVc5NOcEs2Ji42/KIZjo
RmYqaCsfS78Sej/DwFjCyq6r6lTfuWluJADwmgLr4cARRvNmrjy8qWHKDCiJC5Dv
4NxVimd0detDEwqipgO2DxyGlIVswLL08wx7bK3Yl5nLTWS5FWGkR1L7cSBeGdFK
XF6TGvW2sntK7PEk/gK2b+usYLjqVRYfHpLH25iNscjtxHo9xiILrbXSE5STQeyB
+UEpVdWQFtKcxrx1BoB53JoNh53cX+iGqszVGQTpo1XQ8m2VYrCLedblHpjCcTd4
isMb3RuDM8kxEYUFYKgIHjJKDF5YyVZ3XW8/4pWPUhT68HfScfOvn0mFR57JWd9S
SXbJguV6zrrgv1wMyqRqn0tvYO2Kzb50vy1o/QzupEnUorapxKKtV0cB+HOxuu98
xnonRMTFfu2vNil0ebJ1E1csWqVNMmv38ZjAvIO2S5JXPHt/U65Z3Tq2JPGIZZJK
ysMNGPb5ajDRd2TB6fw54kcAqUW0MdHXzi/DFfp8P9rtqDx1iaj4xD+Fsq4o17ag
bJFQLg1b6wfXcfRRc0kxhnvtREeluW1lBrG3wTV6JvbTDTvWnA7zT5+eeD6B7MoL
Gc7EBNkTyPHTjjrnBlllD5ksaZFBf/XtavpDul28smhdmkju0AD/nnQHIlWTG2C7
FcqZNwEwMJfG3H6GX84xtyk4JfgYSoYb58UXyJTj3U8CCMqPWfL5Z9rWwE1cYxij
mET+BvHmHq8BDe85f9azwP1aDa8EUWyKVfR1plqPjHNqqWz7/O+TXAXLD5encH2c
b6tcQM7JKhpnTMZep6DYnOjSXrNoqqtQVGmgDhfl0fcZSU892Zs2mtuew9dPVw7P
Cs8G0Xdxy4g+DroBPGfZoB5SGU9LPW7W56WvJtzj8xpS3MTCjUZw3yy3b+Isnk5B
gmrnIZQFQj65qPnj2TCoMHE19wsR8WIhQ73KaLpXcXTOvGnOW5UfTwqEpherCoii
SCP9TCz9kUqXSszvYO+RV6TRo8KC/ne9SLELLITKL5XYRMSmjeSz73x9AJztBaHJ
snWgyRaHQTjVu5qL84EcUPhWSC6lOcfJ1c7OyBXZYetXJodwRpF1AHD7ueMrVYEf
Pkz2o/+kbliwzOX9w53432GF4rzaKZsl645ceLD946LFcZQILhTJjiY9sQI17INB
B/Mcr3NrVscCjM0gkN/x3IKJuVDHfoBs7ghl5RtJyPitF8ZuKBX//b8g35dH4sBB
TFxdaxp5o5YNf/DSQQvXgrAHD1aYefgZGcJ9kxaXMrkvZDC0ZmNlB1et4yrodOR3
RtDqnHv7qcRBLPDMdTFbmgkL9S06s5MwQWKam4CbzM8LXtIOxfxPXs/JO/HecxBL
8aVSS3FP2itCvVieZDWRGUcbVrk9lrIDZxcDNDZCNhcmXZy8RXX/FYGN6ufBSUzz
SaXzBF1cTAxK3npO6o/4jbqdZc4LGXPsiNxUSiUYg3IQT+xNIVRtiM5CfSvlUz0E
486g9sXakXi5du+BnHLmFwpS4X9CKcKgMc31vsHu4XalySGPXpTI6QmORyAYBLXS
tiV+cTljhTvvUVS8amZ9eRSPosECz/8aB7HTqblX8vWll4HjBG2ujhdPsNLlJv5f
x3UHolkNt8Tr2RM0Rv17W5yXnugsIsfiIsQyggCU/CqZUigHuCfqyW2Ko+dcsi5N
GdR+UegI0BsimIZh+Oxe3p0HsH8IXpSyaUtmdhXc05vqYMIyWVS2AnIVE2AItJbe
Gs1OgMz6D8bIdJ6vo58wnjcKBAQzQTLvh6+wZNpgK7l78qEcrpPnpiydROwAkjMk
uQ9JdUMBovsRXtAXNxPVRI+NeG25bl1OfqQ2ilLyyWFepy9L53mLZ9e4IwEAGUqO
hL+yrHCb8KmxgM3oxmfiTmExgyuo6wIDo/Nvs72Kpuy0V5M4YD2QqtfyO1B74k1E
PJwx2hoZ/XdRv/CEbY1RMZyscH30gLABFc5i8w8ZSbuG81due2gIRn+SMAZHi22G
Vm55vEvpRx19zpO2jUA49ekDeHMzTK2QKJXh0pRXvPAsn9BHCh64jbpfTLyvzrOF
a0LH9Rl5wzYDXq/NTu/dRT1VRrGYkVPKId0CQ/Xcy7zpBioH/+YU5y7vOG1b6IoR
bLEs2Vqn6AedBCo/GycnBFNVrVx1vTdzfqCop20MdZjvhp09f+uY82thge0JvaIg
9KsAL3rmGM9mv/STOmgXCMItNbohpmOPRqaoUWDXjjY+rR1HoKKo1sOA3HrSOMoP
aaSQBr8iYZix1W0Z4bXVLz6KshAgASthTuUe4jygPxlwUGfLYzhihcEvB29RmKUX
PpL4rhYRV8Qd0pz46fmC3ksjLWzeD3rrWygLtAYLn9f0W/wZezm1vynDwn0iKTwQ
SCZPZDSrgq1WPPL/ro5e5LI7Sa/FNKO7/MViNwhNg9tXdlakH8fNIj/0yV8bo8TX
nI+gNapH5oqE7IqppRFdKDqp3AJKS6+dbqugqtPMmuf4KhFKSv0quFEj8iAc1ACR
QKp1BXxWc6u37v75kVQZbqAiZtSsEP0CVz0Xroohpa3OqpVnwoCysTKPP+wBDQEX
Jf8Emy8NTvknuM4BZqi/V4OFzXUZV1EwnZpENNwR/hJLqFO6aSfdPmbe2rKmClu+
wXjCXcm1QmUr8IiWzPmTFA46JxVzKxZ+q3e/kdmK4Mfp4o6o2EY+h5vWKKQAsMF0
m5LX7XL2cwBf+7ZFBmP4rk0eyDHm2015a7nrkoY/eUS/cwI3eOCo1XG/uq7Jjixi
Fb4dAYvlfb94GOcYK9Pfhwop8qVZ9zJiCL90MCU6LADBI/aY4T3jBD1LW1c3Pnbh
w8yQhRpRt0bioa8/yvjyZ3zPYZSZ53HiSI444msORcsY/ytetRJ9l7hKCFdBpqwL
cAN7g8aYUf8VvjoOqIRYMjId/Bg3E9cCJZn6lSu2sCzRvv9jeVvN4CPH0APSYypo
pKxQZ3dJPAr3Bk6l/kazi2TFfvo4TogeQWETQoFbKsuw/z3rccm3s9Pxy9Tcg5Tl
kb0/fvFA69yHc7PjdjkRC7aW80PbUcnQlo6IJ0dtSG0ItESYZHw7oa4doPM+THTO
hOeZZVMUlRhUwqAjk6TH6Zg9hUA71+0VQ2DExJZUpGBPIguJ5/QluM2D95A8y4j0
GGqO61fuUFgu++ZtlBMhoA==
`pragma protect end_protected

// Copyright (C) 2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std
// ALTERA_TIMESTAMP:Thu Sep 13 06:32:39 PDT 2018
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
A2SdAVLgOpT8lHhhAHrvLhKB4WUfPMfy5asGfSBXXk51hcU2OXPWDlYP0LjddVJW
+8UUv8Z3UhmZoiLkXP7VDtTmP9hO0SMhM38eePof/xPJoZd/I9EiMmghTtpslFp8
y7O+CfT40H4A6ouNDOPkPg85xyAOBZ2UrmHkrzue8PM=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 7088)
weak12Gt0x2gHWidDducupde6G5MOojBW0bocV1PbPkU56cXsRABH2YFZ2y+XexT
N8MKFactLQ0TzOQWFe8Dv03eON9TmtN6uY+4kedakcHhvg3IDbLUUMUFUjLTtk7k
s46nWFVQqI+Yb8aqi2Kat3DjA0BJEeRLgVSz5WOOhWFKa5RfYY3uNIkagoa/G96j
e+oC7dhMvhSroM1mjpT7J9bFQM6wsUzRKA9nzkD1UU4ky9YFD8lfl5TKOAtG+X1C
g1Vms7RkyhlC5/SngtiTTe7nHjUlzyI8lxCF1ghysowER8r3lqIsurumdLVW3nl4
XiTGYgJCwOCvKQusxYXvh0iNT9/4/ICU3MnZlPCa1Luntf1N+OLEULkiFAHGAJo7
LO2qFBUvcZdtOUDy0BbDUyJmoclm7sAPRQWdNNrCwK/jJOrtZb7y3In6hiZjtiE0
/EKyAvIU5kcD9JUSS0hdYj9HjBvwYARkDWl/yJLHMOTfF3th3zq0kFNweih1jEdG
TnGbbIIDVbkA3Fvcq9eIvBN2w0+DZbthGPEhov7whAnZ5Tv/eEA0MKAl3HFo3Z6n
/wVQZw0vz3SXAMVAtVdgsio5y5IDa5LVJgha5Ii9ATYnF9yIqSnSR4Wrt2cyaDN8
UUC4qgVfnKvcB6kWAOoGwcjwEUqs1RPZP4wSSD/KGtFgHUeoTesaGaxWyLzYljDp
9v7oLSTaqjWy526cJl+5UHz2+soM4OxTcsWqOBZ2B0ZlzlFc6S7lJyCCbPPhN2nu
SFZKQLF1Da8ltfUUWkn0ZymB8uUv3cN0XmcO6bxNbDIBaQDDP+K3O1Q4k1q/G0Uo
b7gpfNFs3JGmmg+9EOHygUkMuPq5W/kMrRs6Iklp2k9GXHGFHjKg8nRcfZRHp4FX
/8Drn44vI+6A2biJl9p+roKHTDhRaAeNazIA51dVlcMgtO4NMhP/0HrlIDxr9qjb
Zw/YsbS9BkXVQ8A7galaECdmWjEiHLy1tqtiI3mmMRP4N+1V6nQ6hfK5VL64ZxCP
lPFEv6O1ST1iOPi3GllxhFYh3f6usfsQcgbEPid2YoSVPqNeKLVTdjIDvCMz5Ryd
qOl7YCMWv2Fs6qwgnOzbiZMW8tSKprbQfeJf54GdnqXurMbwUe3ygE6KTgoUAoGr
A30mO785UW1gMcw8d1oBs3HCeDhSIDVBAGn629b7fCnk1VMIuQhI1ZTS89kfaR7E
44XiSXvk6k+uugoWIxGfrvNMBgE1KZFfKeZmyu/DKb2UT1vOdqU9jjc36TX+gP1n
biPwXlLBzjM4R4k7cQuL0UdFghwiHINS5NW/ZugJNGAxcttBNIA1ylpepp410Q3F
GDCMRCBUen4t/fSJzJHUeJjDxpowqizUa5xo0QhCQMj15BSgtK/LGfdNIZoDR5U1
GUpV1sexnZAyj7Ch84Cm4KDobxdjct9zyxoBlBjYwUtIK0Hw7FxMOl3HwprE4kTF
jsqHGl96vp49vNzFZ2kvGoQ7QFOv/AXXSBOECHL0ZETvvpAlLlzjxIz3NIZdXDGw
KMZcxbvBuTx746A+qmL5N3fCS7UE2KTihceOAWVHo0T8aedRORvwXKgoqzUVeZ+1
j/lQg5iy9Mi5IjkkCeuLDxuH5cwTa2OAUKEDnHXtpkLd5UgIVHIgk2LABv/qMepY
HxvlksRm/3H0QGqqupz8VsAb8YCEsMXnSGthyXh9HZCV77sqcWziY49NNAycb8qe
kD71ulW7DbNgun7H0p2Kh+unUQRLg5GD+J5tAz8tKnW1q6N/eQNwzoWWKQkwna3E
oa2ZCJsSsOLTYMf2xyv7mX6fgNvcwf+ZLQOJmGdNDGaXLMX1mW4Kx+5f0p7OsoAt
hbOeNBO1r4CIzJEUytnVdtiXq05lYXiIofq6vk8lO777jdaJuv9wsUFnOWXcxCm/
Ec8wBc6Zp/bnZQQZCWW8zwJMpOcm8mqSgNh0vPSPmOkuYwX4pm8BmSEIWM3SedY1
5+yqDH+3ba20DPhUCgnSXt7SB3qzCcFLNjVhrRJaEJlOrMqzj9FuqY72ruFiyT57
V3mWzmEIds+FGF30/FMk7PhgtbOzOD/qiboory3aoFZdTxMtJFkjytQX8Q+Bte3S
7abI2NH2Tz62eoZE1E15YcA47jkUToQHTMU0ym3GwkBXbf2iw0bvFd3AEeB+kKCv
4jERELWeCtxugpGDBzQw+Ra9JySmC9/5qIXZdND42iowMVOXMnZJpQWOL4f8m2FD
dXoZp05outAsmMN+UmqYVJ6R+aUb88TVvYdGzCs3W07fbTU+1NI5uVFbvsgUXwTk
cRGS5cK34hBKS/qyrPKVAbGwoW+hc7R07JIQXe1avc12YEBv1ork4dlicfyYncPu
2fLFWcgRBFfo/lNxFxovlnSoxfpAPIqFnN3Wal4P6cx0vG14m0ZD2+l4x1Y6MtM1
KwXKp0L1yyvUfimDdIqP0yF5yCn0upwaOcY+U7hnZr0jUCD8gTlk/IkDbkBZv+SO
xjmTjx4u0fUVobvihLK4SFJ4DmNTaBauVZnIf+hreheZduuXPZtu7fTKvVJLqwWp
x4dTEj/tyrSR8HVpLyVBQn2FPe+UwjICRgzmErS+mbOv/rA2Qw5/j1OKD13/DI6p
CiTbrB7ADYmsp/XiK0X8UMVHLYFjN3juVa2lndzCRxfmriIusIyO1QimkDHuhiDV
89mh1lKPEy4Q3Nfaki8UUS0lhCBN0mXfW/dvHyJEYbQqSUNHKnHnan34jcs0eebm
WXQ+YAfhS9a/B2CwW9HxBJLLo6XYm5Imrewvg5931Rzrby/9lnXRalfSMFiIr3Nr
ZQDctCV6fWisMpeHTgkLbbFskVFuDd19i/OVl3/EhZ+pX68UheKvYhC4McB+hpmP
mwbYxlufEa3i11p9tW5V5SJ888vw+yZeVw0g57DTWSkd5WNp+ZL7bObg+eSmj67e
DBVE6DMVLoFeLLK6hvRrohIZLDf49M01rr3oqUTDLowoQNSjkNWXpS3pyUFWQb8H
Bj4CJXZYzpDAmOgDiQ7Ef5EdN5/HU3/8h+JHrYPGO+XKxdIROZc7Mb63MjKEDZys
HO6mNllb/SFjY5flcGM49B2wdAILrSHjKRZ71j7dUTQ87UUobAQX1k0Rs4tVt8VZ
5IVgr3hPOHyuMShzqqK53w6VxZ8HK+nUwW3qjEX07ypKaIyQywQ9aCn19rsxBxCL
4oEZJPsDxM8c80hDXkBfbjV/xyQGmaFQaMlsfCFhpbEl3fcis7EpeTMTFAyD98MT
PAaCSJdfrWop7lz12v5miKNleSb0YTiSH9lL6ry0q5c3u9fwx2VlwheveXwexjuY
nWtvhNFTb7fQ6qYhqg1f6PXrlXZQYIzgINNlTifYC4OS6fOtlSKFhDIHUt1nSR2/
bW0j0Z7HDrlJW7EKo7md4UBg5T7dNZhK/3Isx5cQZj7joFOviME5uqkhv3Wd7oO2
uxwO74J7Xe7/5hD6JgjRZNpNMgQo9aNuPWjhkSTKnOAwDZR9JSeISRkJRPq+T2F5
VCJ6acqomsJhx6/1mmmIMwkIpn2uJ9GxOVZAz3TIZliNlBJ2vMFaG72dKnkrstkb
l2RipAUqSf0/xBCWakxPdxqxpx/9+XmzoOG/fXolekCfspCxXT/f679dn/kMw4kp
qI//uaWagWn+yXflmIraCZV73a0taxY2XCMaQZg2LZnG2EUiuT3flUhT12V5Au5g
+zhM7Km3wGQoA35r3RFvp1ECGtapMjkw+j2/Znj/BtWj2T92WRptDGm+FFT58DQn
07faSLzlOGe8tNQgOxwJ8G2b1wLVu/bj44tzSK6qKwOBajAyCCRcPcDXO3OdwGWB
qAhHejDYOik3jT9ffiAwy6UHz5qddee0uHI06O3wHoyFTOzbL8pJRiQ6ocMWH4X/
heVus/7RthSJ02kqZ6SBqKQtoNiJjDSby9f8Ont4FIJWrHxtMbyS3E+nAW/n8/98
0a1+Y0Dr0FTB2S+vhgdRGzEcPtBMHyFfJ4yXDcERpdRgKxD02UGvcHl9j4gbQzbc
wnS4Oa06IGpa13f9xLSNPJ+jRmwVdbs+AYe0F/2NRMhJuV+g5nbSj97hVuWM+CDf
wMaBAzxRIIJyS4HJU89Sk348GtdsIDtSwZ5LaMsWkvuodfn/HCOGqv+wWFwzHUZs
AyoUNziRy/LizC5ohaCaZuYUUMDhdXTGeaOfHxKA1j9yhy6eAcSf1t+wCDYfI2PS
3jnqIaNmBfNgrhf+QbmMhWQg4+Fw/g9jH3ik9YCFQ57UHn087V+L7Co97qKmk398
Rps1576A7zuq9zNjtEFCsbEgwUStrYqelioeCJiAoWWNI/5rt3KiW/2SoajG0Qq9
5TjDCdwZUG1NaE/vfingi573lS80Qq6QXw6uZ0sAyLVuPGaiReFrLj/5yZmHfOhU
T+QYeQnpN1Tz5Cu6OCPK36d4/JHEnO73cvY+JOh31fFtif4ia1bZgSF2T4c2SqdG
tXsjk+Cd0yE9zJYdV0SSl6bKyyNaWmNeCA5FxscYiYe6EnHu8PCrJ2OsFG/cCsIb
X1lF1Ybk57yM6j6OKou125ZDhRZmhjUDL59pdvsHrzpF+tfdm/tG/6ih3vOSWhOY
jHWdNJfkvUWXJF25affpWdyZ40uHkHlJkFDGffS4m4O++fE7KiqPx1IfwPnyzHni
sTDL3mMKmW/q7LtwWv8jcdVdc0gaZ4xHWvkPXFpHp+iYuMGfKk1YBSYcYdrRDPpj
fB6L+svry/vE0I0R7XCNXesGKsCGPPuFvvm6tleNKaWsf9pkup5JvfYwh6kiF6hb
eZDuoUs8IRLYYOKg2XGc+kg3TnCSDfKm6A+2pYsteRzuaJ2C0qBvXkDtUVykywTb
4sIcwj3cbn2MzX+1BUp2UCAF5VwssUUsKAL2UbDu+xvHv4iZXtkZKzkP0gFW5AFm
6DFYLI/M//YabABYb1DI4+JHuzr74xDVpkGOMti3m9Z/FDOOZj34o5I75T082TN0
1/mrRwJxxHaq4xfg8o8jT4CAICkhpfDYAUYoIyMNggPARyzhoDI4exni74lYyNt6
Vu1iaOyGCkKDYTmXUEPUGXRyWACtzuMuJ8Dncrrvybf1ohO7MksF4xz515gPIwj4
trKfmPqKOlwPQEaESvDEPh3S9laP+PzdSvyQ8GqkrJex9kEgd3vDqJJ8n6JBU2vS
ucbH/rI6bnn7hbPgxoTINuFjjzzhILb1YrB0grw8YEVEh1gI/EYhDfIwBM0550D2
iqNJb8fZKnLosVOLeeY4dK+H4Z5ge5iGeH/QTGR7vLb/bm0RA0uRTObs1OvGQQz+
u/YsbIbJA+qta7kzw2kORhXbeLDkU1ux4IeOp8wgw8ZeHjPjMsEqP/zF2fB3jvqe
Br7IZlPbfAUuAHRBb8juKxjanNm8RmBlzDQs1uHKmoFUl4dhHz5Rk/7PtO4nc45F
r0nKN22H2m0ZU/AZLvuB21u8fIuRAuBW30P6nZlr/eZvkzHcMQTgHAXs3SVYlUFA
0Y3FFMbjS/jaxA4kHpaeNYA6112taOTcEhOntXDqfAbDjQkEZN3yxmuPRW9rV5Dv
/BXjFpOpR9v1n27uMezkX77abboI+4BnJByyBWgtZAXelo5GPDfiu1juy+UUsywQ
ZLbPUyF1Cf3AFUGCvItQOqAKPWHvRvjFPf1WFjLrE51OXzEfftqBsRDQo25Igqz/
wvc2wBoMEBQief5A+6cHzjZNO6MMKoQ+nW+rSlzDrGebXL03TwJ7/m1wPghr7/t5
k9HF1d9QM5G4EhVkp5kfZtNmHkXtSh3Ybu9jDuBhUpTXW0B0aZerD6NVYqht+6Ji
UZc53vkSXom8yUEISFyFtDScVhFpsrU7JEJPyGrtQI1jL/VVjuN5/2nRAispuOuJ
HNvm7JiuctumG8a5dPNh+IyIjszViLAAc1tK+fDEyAnnWD24+1lieHqPuDTC8AOH
9od1vLsxK8M8bLP6tGkI1s9oCavktdEXPVu9xem8xY7EkRuWiii8tm5uthrsywGq
EWMPAi/HLB9ev+W6hCeTtAe0iSz9rGBIbnWvcfCT2yac+rgI7eQTOUaF8bouVTY1
Rqp4VzW1zIoX7Ho6D5OWrRPSsrvaYNt/dhdIgQElOa6217VMljg+u5P325vqn+Df
FVckHtmY6VTh+Tt8oem5kNacLgv1/Eu584oYghkx3tH9bEpJQRTx260ymt3Cimto
MrhDLknxSbmgef2yVDYmjXIrCBeSDfvju864nGRIqr449kQ8NqDC7GSKLmVonAqP
4cMBiekO1NjtW4KEJqrbsLNwUyKp/OVuz5qZBnZXP8EIp1d1b3ggBiM5nmphweud
ikVZtjCC9C5WTCRtci3hFHN9io9lbeWkkqGOIXaiKZTcrtrTVQnB1qxS8Y9WWI6S
/HOFEbspQxtojve9qSsh83D9UXLUnAdVQCSsDn3yVIIJb146qobEWlS+1utS7LAl
1a6VZSwWZGf+b2PIcVkrhjSyNdxJJmR2oSuuVIXzvapREqpFgNNEM9i+H3PEGa9O
8JNtVQcXXK6WIti3mCcqsh07ZbgshAg47NO2dxhqwvmipPaFaPTPEMUXKyMizyMP
SLcr/n+rd/wXDFNEJxiR4v3NB2vae3t6Gw+f57Qyr4oAW6a2tP0YNW3YE73c9yLM
E8WD0Svc2cD3L2xPFaHUqcTUkW6xp7QAmnPdfuxEEiHp+qQxyDDUKqNuyCgb7yB8
EjzjsD8UEdhZetsHFqKvn9YFQq0lmq6qaUWLWUs+snXTdDOGwMHxqtMQHT70dybd
ldg6DFtPBCl3WBQQ0KScfhUwixa/0xfxgJ0NYUz5bkrQlzJeq2MOa8fhDmmsln3P
6QvvSodVe2AqmqbXl7Ij9LdGrMbL5SxzzZBrAT2Bc2bCmXJkpH9QkmoB0tQGZwzY
sgbal7Gmm2SlUjNINKA/dd344F0NcCpq0tLikB0tg+8fmeP4bD/vRVHej2996/yU
E+lEB6vwCTgBjPneTMRNTdcuvh4OTZXGhttm/lJpN/sTO+hmIsDlWdpbUcMnw1Ut
TnuATKAF3GJf1YxOerthc+bRSdnvdMFBMZAWWXE2TAYil3IRaxcYXOKBKD307Qln
tlBDfPmv86/wOuoYZbpvwZmD6Jq52SlkDEkaFs7l8hmv7U5MF5qh+X55u9911orA
VRKVdZOnYpGslkie7hD71hlzzxxbpYdXdyNBJ2occ7+FwQlVoVxt7eudE49+KU7V
gkP/EeYjMXjd4Ej2vcFRN2V+8YtjKMzVPMUysPJQMpE3clZpbcQ0buBUSmQeFuqc
deBpqfNccpza8wCAS2BQR1HbvxISsz+/NOs4JGc8akQYQZ++p0QRQ6sjk9ZI5xUc
Z2KYVyt6oLT2gVqGysW8MWQO1OPJMK7Hi+BOpZ34Xg/RF97BN8Ny2n1QsCtYvZjc
X9MfyTS3ee+pG9nXCux5XPU9cwvPTp1w2z56D0nrJxHfus1WGlMyXcvP8psrjEqu
YcuunvCqy9TB6bm9dBY7SGVQsgE3znNPPOgxEhJ7A/CjaV7i+XAXTWsV9Sp3GcsT
RW24zUWcAX1GgohNnCS1vqCUNen9HB5s+EXjCsWifHUxJirSuqoytOpkuTiSeaRW
hfMJJrb4QRp+aW4cO1aKwZrb+8HLkegOlTW0aCacaCZ+RopOp2YSmUho50DD+hjg
aibnxfUTT04nMkmMByvx52qL1t2xDQY6Fs10K9N2JmH9c046vC2K7YSKMsBpB7kS
fHX/CfMiXUJkeCvn5b596asNq4HYxutld7gsVcl0q/zw0M8lYoUcOhOWWk7DxNuK
nxUKChL5VggSTLVNzRhAmH75eHisHnukKlVjPGHQj6JHekIRZHoHwlg/auTNjTSB
qryPp5OuV9gDPShrNm+xwaE1YPp34c77F/0kNnZ6ruP1+9w21WZjq50JzIzG8L41
C4VjZFPXq6SWwATFsjniVh3dObUUdbDyP7VJpHgXJWSZlqW9nbzgHpqiEmdVwm4O
zmB0DBQIRTEuc9p+RCWx8WrjiLDeqWI9SnVKjiqIwKrgvRXKSzluNQdGFMdESTuM
pfIbDiKvbv/iFCIQPFu/1L8CP4XiXijRSjpZT9Ulf9FWYUEq4yfi0k5McENS+0Y7
0gokv16zGlHhAjbb+Ll4l8ASyLz34hGM5XxYbSMw5frf4EZYyducHtKbKhR2rVhr
SJgqdpIH8wglm3hn7OkR0vnYcFOTUSsDKlSqcCNZq6+t0CVRefqmFzye26PGa76H
bW9/cpeea2qmuTGK0UjMw5afJv0zRvqp8XdDfGyvDEaMT3E6jTKmby8fhUJyY7/p
Ojg76p7GsUDJ4w+UVw31DhKdTGG0d29C/5zRMCdW78+pvjsH6GeEynDjIVHU+6a6
m1l565stYn+o/vfC8HK/EH0auogOc5gc80Ih/++hj7/viMVR4rgmuG603JP//RZY
kZC0GcYtHatzeioNrZgiGN7VMsI/1FwjcJM/Lgnq/SigN3vtQpTGswi6GNuj7/hj
0Wmezv0cOZvI4dsog9aDLiYZckRJmfnErRN1AdljAiMM8nxoflK8qTeCtFkNTAbP
4/YH/SGnfagLa/4sX7PQl+fEju9UZd67WVTOymLk+4LdizpQyfmbdaY+0gzP446V
lyelT6nJkEhe+R59cHeNNX0vkcJ/crSVQJ71txVSR44YNpARUNs7JlXbSXXbZzNP
hUCdEBZHzpJEPIod4ybWWTIeD9GdHp20dm7D2GLBFjzLcwkRTNSx5KXrP44N35Bn
uOVz2I1ubP5FO1TO1O+SVYd25vlkcmuOCbrAS22JEpmRDx7dP15rsSg1aK9Www4j
GFQUPSLfSolgcXShF1nvQ2+B+BIb3t+28/WfxOdYmLHIqoe2fGFtxtpYzZ6EXs32
VqvLB9+Zo1pFTOQ1ZmiJ3IRU7LsxWFtqM7rDFsPNkYpZQFuKVkUM1XtQEtDxgKGx
33svtX+noqC8auW15XKo7mllOZlPUImtetpFD0Agb4z1cqnG17ReAqeaUUGwE1ql
yIkg753BkTBQhBahcaDZvZh2IXWokKbjvqURansuj1X0mb1kUAmmB+cX8QAHwPZ+
j02Kov1lmfODsuOc7Nq8LcNKD/4vaQawgzijhwyRTjqLTrTm/7LawiA091lpmhGr
WyiNEpOp2++IlA6IQl46PYRRbW17jEQk0+2XWjl14zhGH4bPSSZPb6VErXtnT89W
+7eIJu5uWI94hh9dtOQr7utnYpmjKcU4Fckmf9HIM6kStrgEELsm4ZMHYSG4ugii
Jg26lEBIgR9sHUz0k2B085Iqhf/fzyU1cYkzW+BhGtxcfPEzaVdRnDU1iGSkaC94
mibLafXO9jJKaWmuw+Sr9oLCL0JZH9LAmhASeeqFeNR5afoPpKjcuOhx92YArQnq
2fBsPsYhnGk3b04wlzBF8YEZDMjs1As9h9IFNCMtlJI=
`pragma protect end_protected

// Copyright (C) 2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std
// ALTERA_TIMESTAMP:Thu Sep 13 06:36:50 PDT 2018
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
PXilGo5Nlx8rijzsHSQco9IHzSPdKGPLmynIS07k3WL+/yy9+LKmKsiDzMqqzExM
Zm9tZWJ2Ezh0wyVpVNnzwoAE7cVaYG3+0HDP6gbIfn607Q3rjRDx5ifGTEd95Tq+
Xx/HC58B0TySOPkUMz+jMpPZWPRWxK6cx8lQIZFZmLE=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 13568)
Nki9gvgOwoLPi7bB0T1u7yfy6NTnSHsAbhGFwS7fepH81pEFcj2RCXvfO5DWWPNG
CtQ+9W/A9BMcNpMXMxmjdLsi3zn8QX52z/jLwiCLjUkQG5uhY5caKLRgDjk3lX4g
T51wiG3BZ3MuBp/hmqwgLiYKTlYIUTJZYUzVszW2Rr0OYN4pflRrtTyN1lU+enuv
4wIQZ2ggSskxgP/JLE3niqZF9ksUpAbM0fFUonLmxUPGxuU4xPHrku/e1ayYMySA
v7Bglwbk1jLiQSTXGDYXIljE+ru226OWDJyp3SiWAZiO5GgdLk1VfVADHY4BHZOj
FXHJemO6urdFcNyvu4WtD6CgeTpln3KlUndCFuK6BCWV5nW7iyvBjMiemUTIc7CU
CG5sY/xwe1IQZAvIADB8maS4y81zh34wB8zSYW+X3m8glCcj8qUSsNyVyOPpOPdE
3CM4Z9bh4y1/zZiW73D+4RwUYwNOfvuwHiIvZTywgvNLManNqXX8dnzZdjhcwjqa
nbE3ObTgZk1KgXt5/MBtoX3HWpOBq6hpyZl+m6cM3TddB5GY6EcVScv7V/psV8wI
FQvx4UtJ/Y0aIbQEyYBN2+dGH9ihEArl4d7C4lUX+FIXm8ra8PKWygwi7OsQE4Z9
Wl3JgPQU4caQysKzMhEZ3J0/n83e2F7L4NgZYo9YUetRepTvy2cxicjUa4yIwjJn
sa5IX1uzf3si0zJ26PuInkY46kkQ0+WZyhn6MSBESBS9flAKgE/GrivqVzYrZlYg
WaC/I7QYJ4Y3yTDwT+wuJ4BuqwyrwJcLZ671gHtHF8vdfSdBkzk0P0WAHjmraVFX
da3CZ5fSnHUO4Btyr0zJC+HfZNrWjzzmwfioadf+DseBckAN6ujV7LC3MGlR8VMK
G7s26BYOai43ik6O1GnGq3fB2Q2Dc/a7MG1z0xLXAFXT76CaZ9m95qDs41DPjTzY
YQlKlSPyIOvtMoi68QgEg0I1TkDm7be25FVBQARLihLhN1NBnV7UBvaVWPJxshUk
MyqWnCZOJT0Z2qFAhrjm0PEmNsS63JTbsKbc8mEmqG1d3EQ/9GX/B55XIc5EtacI
25g+Ye4ag9zI1oZQCjKJ83/tYCgYX5Ym1hO5J6Aj+YhbECvEwqkLUBAuyoRvI3Fn
z8zw6MyijK97V1BAkpoDFlvjDQhbL3efOs6F76migbgT6wISiUC6SK09BERQKqgF
2x3CtjhOjZgveNxax4iSQq9bYqbtj+EwhIs4z/xanlz9Eke5gi8CTg1IYelxvp92
sZiT3ZWXBXsSaxARN+db7Z6cfrcn1bVlXHlTwIXr9+Y1fq1l5/UDCXr9oFI7Xo2R
Kt47UEXPHdGJ4yHBPIHUfQCeZPCXc74/QRChCmYk8acE1jgfvBvBFR8rEqsUhLwy
sLrTrMpNef2E+AVksfQKRuIoyRzPpH+Stqk9uSMT6LGICu9Z8++jrmzPhODeLbSE
JBiViZWfRX0ZFriGMa3JQnP291yxBmTNBvudclq132YEkv0SAt0aEtsp+oBUv2WS
EICNnfDu7FGLJq9eerl7Fnx31kt89aA8RYjTYtwRO0+3mhSlVx979jnAWoemCSfj
3Isg3gsQG+VoHnTHCzlmidG9pooJp9KKto2/CrfwiYGMYYn67gJgKf6cD1Y+mBaw
g4v6hgaIC7nsr+NEg49cn7AWFLPdcgWMXsHR9IcKgief4BPgrdLcXcesBIWPal+j
ZcQf5Yw+RoA9iGLsHGR7HWt+fUko74JIyEN/AH5MoFWn1MEGBnRwDIKo4Q4PaadV
EcDZNIwCAWH2PPhl4CgW7Bj5XSQYPr5vQ3y8VWlkiKtFqf0OZZ2DxiD/EZU0+Lpd
fjHESoSwCO2DwHflYEVc+r/piHqMF4qFqfgjIeMdFW9aXpBuONXULhTp3/XZOmLQ
EQ+Wiea/pktULLE8mNJFz4pL0rxdASBsjS/ejtx05A9t3icwh7zCO1xWro6kCOuO
8oM64rPqRzTxn96qM69m8W5AtSfCFNGQuhHjyaBUcF0sySzUhHmTZ4ouIwNsxCJf
JAZHnZlmQFjbPdjwL7uZaWeeNrXw2c8LalbeR0mTiugJb3aIFiqPv9+gJtIVIpAF
LsAKVOwdC5xtWiFMGhkglh9t2Yp1oxIBj3O1IE9lvPW1JwVtoNrg75bZRK8IcXcb
fPk2CS15OTKF8vcdatfBBkWKJJsTje7c1RuAUWOvkX8CF3KmFC6DLofx7gtBjc2A
TpZkZVpCJasFM4NPpntvSF5Fyz4xeXqlRDtCD2yIf7Ys87lgUjXh7LLeHBoqJZc9
zQaLzvOiivue1aqDikSu/Z/9XTWOQMjj18uoaHF4t6cc2VX0zKQ0J5TcMkhbwC+b
K0tjrr+EyJ0mVreTmJV6k9zO6VY25YXfRTKhuCsIpqXabJSEDOG2UxMk6bqCqBgI
wZldMRa9sG9oBqwHBLPz1Voien39BrdcznPXRjmC4PvLRVx8O5CmvZ3aSOM+2sDk
EpcQpljVg2SHARUuVLKa47ze9tdO7GxF1zpnaFYQGjj/qn6QSgfBTKYa6YzWNIqj
EvG8C1rmNhU5mrk/vaBXxCtH8GqXPQ0KFMdA4TuFSjtG2URlfho3HBwBsGt+nZnV
MgNEyHQeW0r+EzX6VE19x39JPMuh1P8QPQa0Dt1wmD4PrPLssemfdKK9sbnujSu5
z0CVugnrCtcuPeYBiQISH0oj/cwPSe4RzJlcR2tz1sNJ6N0DnhBU4PMxbLz7+4YD
xIhUOh0kOX46+xUzFAL9qV1KvDv9mInYNot6kwPi0bdEtmPXOzWRI+Yr1o3MS7X+
UyVTxuNCr/VNJmOk5/s9nf9f4YRYrRpfwxWBPvLsd8CXYZSR6lN4kKdO/zOcDS2j
EOjvWN90tWot9eHmqm+TWV/H/sgG/XEXWrOcZylj7DQoDx70ApYWJB3FZ+5AJkyi
86UjJyJaigaH5Y9GuY7XDE09E9WWrA8nYjmt6HPDMaICf4y5m1IgHvE2ex3QrlBF
aLgQm6sMkBuXpOPyYtwbca5gi5+s42RuCaK2EC7QdlrwPY+0pLehGVOZMO47wOb1
cYgQ3k2JtPfJp+J0yyHnnVogaYeu8H9hjdmtd2vIecDJUxRq4fzcCh9Y1PaVy07b
aeuxIhdxSPDd+rWrX4SsJ4fAaQ2vzhpkDd5YmrhbuMTqw2MvD+4wRH8Ua4llm0Wr
SYshAzxLlvq0U7ktd7Fa11Df6yvkXJwrEni9nlYD828LDz3ArNSAKLDKzQx3cD5v
4lkva5gFMRBEDYlPPoYm9lxua4qbOYsKRTRvdYka5EWAs/U4wi3bAeL9tIuY20PS
Wr87oFFOELwyPwkgZo/0qXhMq4BC5386f6hg+Fuh4yB1ehBJPgrF+U5rFDcynD/V
1VT58JRxLYcootzwUy7y/ugI2YYaPfBrp0F3h3G0q/0UgSjVgZDX8Gzu2Yi0yIFZ
kXRBq9868JyC9uT+sGgxh3Kk405OOCrjptMjWrv5ZVT29xO4qyG+HaqotnwiehwO
eg9uW7R1bQJA/jjf1PO/vdHxxGHhiMoSRgormWjqsVOT4pGBE0ZiaK0Z2VV9CpvQ
vS3TtnIpbQtkzYFO+IlTE/w37XvNem5KhaitXHo4J4iyKn71bkZRY1PiTYZU5rw5
+hcBZWap7SeeI2PyqYyMqlkx/k4/yh5PcZz4opqo6hOWbRPlRe7f94crGMq18+m5
fQKPjP11G+9rmQiIL6YYPx5bePDvYk/ygskXpKRDRzZxxoAA3V4STAHdB2uxIf58
CGqIkfjEKFGMwWVOHV8D/q7KhWxi7/GEFu6EG519fbmRl17Iv7Sq7FPgvT71FShi
mCetpEBSwOyPECJ8IEKVBhdoxX4vykzf4gYv273WcmTHQGsxsX0IkmyCCh+v5Gwg
OuNppXfmljIH39sZCJBKFo0Gtc9n/+Wd5xvbG0EKut8uy5UNoYDP2PhgtQqhdvWu
L1/4AtsEpGpYEWXksVMBGhNAGw8lHXKwQ8fPHPNrhl7K4Ql4fRHi/E4MUpoEvDEe
RxFIHwvGqjxlISST63oToSkqeJ0RWvgx7oBwY3bNf9TafvJuo9tArsvREF0k2bML
AH7s/6rKHVZkxZXXLtN41nC1NqJbLPMqUqRs1VK95WkkZjMDXDeHdZObUEtYbPQs
iKipaOBHJt9Fk0mY+QWc96GK2yr0KWs3UlHyR1nBJeDdoKBC++9wgHjaGixxj37g
5fbQpxXvXI2TP4WfYouu6kWyiHrVDTxY4CmrWqVboIm/GZU3up/oFwhB0AAhDP78
CVwn1i94KkKaYBPMSzndCA2iR2JN4+2ry6h1bQ11TCmezYCOvHXXf5BMqirhGMm7
wLpTX7YKjo8SUVnzXbf8144580P8Lu4Rzrou/EJPI/hIlCO8LQB6DUutd3HEu6d9
bqOhGXjjmTWJ9tnr2ZENsJ+rvz6XdZNP9JxuJRnFJ4NyWaATF+E7mU/RccpdV+s1
qVK45dzkBLJr+xxE8rC9H8t+zXOZvgh8gEUayGUZ7DX0bxD5U3GXXiQeoXscPyKr
Dxi2kh2R2vsj2OHoFOi4WlwWbfghSHPBcoW21n5ifHN5JoXaUjazw0+/aAFYenOf
QhIxE8dpsZrjPgrBfsRcXfqNTIM0oC7Sq0557LpA+syANDBm6G0ZDgDVs7jRyIMY
bka5rH8VnVcQIUBZ3QJYDnyU/K8A4+/1hCcGkzMxsmpjmKoWrN7kljFCBC8UOycV
juS1Y0nS/07uYim3OOaMP+8pQKYsS34JFEHRJjepTVWxqfcfG+ycFyZaaHpgahB7
zSKINnq0dEe+8U5jH8IX4nxuJLIj+YMib2/pWibFyX73To4/3jGap3EW2gu30U0P
w+ZaMR8l+kXCozgedXVEjkw7ymeMyVtGaDJVk7kaqW1v/zd0/Jy5I7iprucDJjwO
irbqLT85rt7gpg7Fhj8z/QIaK28XwlndcqOa6lb7FPnRfJjz/tY2Tn3F3Vfxr5gw
T+39xd8/WuJAB1dphaWX1M/klkciwzpGm03ZOA82m1Kls12pclFDAFyBRfcychA6
WBEZntT6IDIq0a3DrBxW51rWy1ECoNc3DhjkEEs3Tpw83EBxx7Le0gAz8j0nhMuU
0bW6JqS5Xo0IWWTkWIJdyOJOP46DfoKy+qe67fM/r86YBOk32f9OxCUYbUhJys/2
ld6cfdEKWnKr9mE/ckpGW0tS5SrezCvmzjveIsNR+buyukSskQ6XbOsj339hbOir
y7TbHurWwfHf1uSMVSGrzsqmiShzv0mzDI2An0x/rZhAJ2E2ApIKy53pXqRK0wl6
YuTk1o1KwoNymXID1/y4T7/2WGwJeTHu+WFgktjAV0jMQLQq7q4DXlXBTSTO7kXx
cekn9y3F6+OtWspm1U/qKsnI96zsNt0ZfFPgISOqVKXBgQps0ZGWhWZ/BVnDnkGr
/i6YK9gNLi8yQS62eYXDJJSprZ0A9/Av4vJcw3G+h05nz5BmtUP3PfzlI1H7xAVV
APEIosjP/wmgXpTJdLZMq8tFYYMCOXAxNEcSP6l012//HKW5+fvUIJ9WN5HtXrC4
HBek08zWbTSvGzqdpe2XeMoAT3VuFYBaHn7/EOEsSzSmSqS0mR8xO6neEB1ed5E9
KwT3S8M7BU8mYucjZDpiCKE4+9hJ//rtckvzqOngeXdlPOy+8nmTuedif0+1kIUN
9oTKw8mMI1dBqJHETSmV6Gmim87eofFPYtNgUEPk2/Z/DmBKXdm7uWVgc/wv/fBp
lj1v8eHFg0/a2J8ObdnOm6JehQH/fNk8PBaa2a5Ot+QvPB0WAEEQzY0N85GsziiU
ZlUku5kZGi7WTtxKk1RUDQwryjxyTdGhUIVqM5lXxx2v+yXU7OfiWzOrMPFUhZt0
o8iQaDBjfEZg+Qr0t5d3YA2kKLRpQriwVt7ofYB2DFeDdYMJQpuEx6jsXPjjzygP
IFapuk5qAarYajp3rl3Om03ELHp7b1NrzSrfydWuW3MWZMPTLixOubPVNwDxEU8n
B1xaIXY/EVC50crQP5cMG+whbQrbYSJfvR26LozkAKmOchUzPGJHb0ATCfSej6QT
BXq68IktN8m/CU2hZgiQ7xEMJ1ah80YzvNqpbPtq8Pirn0lBr9U+LPWoa1r5C01P
ly8NuDFajXw0eTcgPq8kZDiBLaEm2XTWNyx2kEeO6SqmSEK8pdJMhW59BL/7puyM
3R/fM36t1n0ukkGGwAJ56kgG3vBhUhzRqLdJvcyfDu13YFesIl66hyVbkckPF58o
1cSVgQqz9TgUr4K+J9x6NULr7jwit/7cmzBYkgNuhoxR4bFx1nVX48FMn0a4NImh
85sz7Ey7zrswYaipV9UpYYz0In/bRwh7kT6W0jMTGIgzejsDSmntLyiFGHaIqGY+
qjIaReDwri8LzucaIgylBJtMKQC8vrlFPiNy41qRPG88HlJFS6z9Y+KHcMkGGVJr
Rt/W/2h82eJeCQ8zfEUL/R4g+GWmU0RpoQfumxoks94+Ppwdmmaz9n2y0u+pSugG
mGOjt1rQbtoGAuXssNi3/86fAAS2jI6l4qVz1w2VIZZIin5JNuSgZh5evJ483QNf
FIy9g78ZMg3QZYvix/TZix/h1KUWnz1qFHkUQgTx5I6Kn6G2+gG+E2oQGXEqrKTA
0vW6hhT7jniXiG0jA52wTuSjFnWwTT0xV9EHhanbSWFrUDVVAjTcu81+8ZIdzQfL
VQD+BgPZHr9sb1cvb6/xlEVeQ8fGbIMbHXurrXiAZR6uO0Nzy4iusyYRVrS5isq0
XwbCljBIDNaXpWToxPNIMkhwZL5py8l8iXL5viWrQQfRxDEgpmifwwsZXULqjvGS
7/77wa/M5yruWe1N2Qg+B+cnuQgnKUSaG7ZTZdLE6Lx41RbgnxjxvrfuC9L7pSa7
6K7+g237dzxTvXfU4Y7TOsyndsdEupyCTOTqlJabmZ4dIcSJGl3/MdpGzlpTcw9s
NDSSUfVWYErcstSGdNJW6rbLHOpgHGTsb91vfrxlakgTPcchRae1ebV77IdATwce
FUiFuzX8lrGmLLIRez9PruDZOfjIsYTc9mJVJFMRMeeXiuysZRe/Y4lclt//CX5X
udmsv8qjT/X+qYvm1i8ig15cpiuSZb5XT8HfQP79asLss8ujZ2hQKenpEH3VauUc
ECkDGDZHgS9GBWJzDAJQYhF4mvCrUulHVHBlLMySmsZ95VOnNEz4+InzJtC7qqMW
rS+RPNCWp38Eho2mcbzTpVTA4IRe5ET94yfu5T+XTHIf6geJmDbpsogAkG+pSnqF
mOz2z7k9GG747YFsas2VHy63KPYhuCAAoyMHi7PVvWKvn5m09ok0JMBa+YT+9I04
vhGw25Mgy/o1WaaHh+5qcOCi3afznbLqHNb7zLfvg8ostua9O/2EXpst0D5nHg4N
+vsOB1HpAlLMDgwH3/DcKNSLVPgcS6XLAke1o5WG2dRNoXJpP/5W0+rww0hbuN+S
GvICtN0/r3AzE+ANrStGHhntChZJYRQRnsBI0hI+4BSsjg6sZcwJVvjBz7uCLuy2
GnwRdFX3IUU884EeU9+8suMBPxqypt/WcUF+bVY9/GgLtEaMybBgyn76b37vEczB
jemlDV7J7pNbdi0TPtIYmtsyvoRuzfQe5nIKebo0fsl3a+0JsKhulzWZ3ggmCqnT
amqcDRKEAzBgLWIHRlAkUdm+movxvQDeQJfz2vNyOzfXnMzgUqsaYBN8FbZMHYsQ
Nk6vJfbxqmk/0DxU9MCE9uEOce1yJrsW8iTIuUpvJq8EnE/LsbmGhrHeP5nCtQnE
uUKMGhhHeEB+DywZVZAtukl5uH9CFnyIIWqe/EzXns5QsuTYFVCa424UUPu/Oxlh
6cCeY+GGvNoiNGEw7whbteiTHYqhAlUOw0VPfsMYq3F5+c7PM0nEkNTi2NSrqCNV
Y77AWJIxZwgwFm2vm1KF6WDtmO6I5lkPS0f2tUTRDsJX+16CbsSEdMDGEJasp0mF
azdGg1wVQUA3HnPn3LyyhIeyjzF0onGBPX08lkb8cWydc5LgR59Jj+ZLnUgFlijN
740hH32jSEkYjbmg0GUVLhsPDglb9KP9vRz7R0epNXk99FrsOPp4Pj8q+m+djiOj
hpPucgv3LWNN7jnaCqSL5fKpwQYqfdTfXQN3qGaG5pN7TO9UNgoyOGUTlEIzrd84
xIS3k8U8EuLvg/J4PSFoQmRID+Do2EvLgktQ9WCSC9kRbhpw9gruNB/AmaDuoQyD
6QHN9XuygikbTRCdOC0J3z1ZNDIdzFOLtHfzJ1WhFA0gkPbsUdwLTjRaUzf09FHU
q5GFcno7K5IlUrLmx6Z9wr9VyjY+28ObukuF/M4bdGdXPyxJuW8jWI/AmJ3GTHCC
2R8SW1F9vI7+3vWvGxZ+rkQS9vUHgFmkglzGAU181fRMEQNS/tqoWBeiRJNwfX9o
/96QGuoBLbiZY+xtANft6bhZGHNnvDikAtrvSPL5v+S0Yt3EVcv4LUH9YxywrvVu
F72hgPpLyFiyqzvzthy6aydGdgripuA5IP53g/qaLQRfNQCe4YpkfBWgt/aMYh50
Y70L5rfGie6Y9/npEnCuWCjcwyKhjNbSWejYEWgQKAF+BjoNNBJZmld2JT0MBZ7U
PO/sysgLxVYoH9UlIXotbTk6VEWZ+b0/ZD+tGqmv5paH8M8vBalvrbU0j4EjI66Y
BSQ6M9OqsgbD5/5SqvbgSEw6BdxhWE+oDKbKK8kiOCO1B0D5pXq2DgALfCnzDamP
GfStcBlg7pY7E02IhSbuvYUZdkqctbT8tK5/2KAr7+s3PewfYEGa9QCWID2RXnLi
EgKNNTgBhLo2tFRwh3Oe5WISbbljQyS8LnUNPmZXJg2v0kRi9uHNKJ0hW/akQ//6
q674eKUVSBA/3E3x/0ZJVi3AdJ2ATNy6DarTSTTfwf7YXSqXSw74l620iM7VqiXo
V1mkqjJJtD2/7MQI+yEg/mqYQ+nFDIt62F7/iAOL4/rK1241lbpwit2XI2yc1FOd
Y9fCeKXzFHmox1Y0qCNCcipzHk9WgfeCx/CY0dTsYLE+pakTBP4VlrYEWF0+pjMT
/KpRi5ZzYtJfl4BMuCg7MHd2dVCJkBnKeMOTZTQ4JWMhrqEKPx/njVRdiet0B6G1
n2H4TF1I2OLDMu9yaUZS/lfgH1dOMoAUkXkBIpH56/k83D9OtCnB/zWMABW5L4x7
hRaQsJXnCia/NJjHxpmEg1HCpTfhxJ/jNo7V9OKV0YMtkSE32qxM2ywVjxVfTXL/
sflWPW1JtMGC7sw1LmdUMi5XJU2nt6AfXlMG1wGyh6zwadZrvskvLy5P5cO6Mnfw
Ln6EBN+/3DGyEbf4pW5V1TEqs/bdy42MLPJdZSOYzeRHI+PSH3UJLdcIgchQqIng
rIhN3cY8g1dsJM5F5q1EY8hm1j1US9LdcJh4tLrP8Gcn/eACU8HNEUJch6fgztBA
CxrwEIXUPAjuzEpor5PWIBF5ivbIWfrSFmxtjz9EG11Bm2Rh0ef0Qe0Op0gBeBWB
4e7vckY6Z8axEn3Rer0hc/k07XlvGCYbSzzkoDQHfCLqGynVzJf4d/cOarZEiAqW
16UmTlXTiblaWgLKTxqFrT5FzlWQ+4hliXvg4lNq8i/wqMes6K/gMzM54hr9SbY0
TIL8hW9/8gKoF6/vSNyaPH58gbZNb22MJR5XgMfFhdQHDwSOvG5HRfPlDytg/Gf6
DXah307uVx8h+7hJvDjwqJPerBOtr1pfHJBg7Bl0my1NKlAedodiyTd/NytdDQQy
B79iBKsavmHSlgqZA4uQLDYvA8JlEP5uhx+2EUO2i8wvI1K7emZMgzU4Ygj/TdHm
So43mXEdw18unuzLESmBQSh0zhkwz4LQFx9hVjKYHYrrbqKoC2XMOxevZSGB24np
WVQ+QRX0e1AcP6jgOxrV4efEOWELbftxOnExQcerIMpATR/fC/lCeYjvjU8PraJZ
2rZ2l/PdQnTwXuGZkUgsZyiERVhdxNQH89wPhS6UoObPtPwuV5jy5nMMWlHDsiSK
Tqch3iroEUkPRk/+qQcTaxaz02s0Eck6DfOCPPU2MknkANtx8yqh8D2xNBNjWUfO
VL8VUM4GAjDwQVded8J3fR5YDeZPNiq3r/Rg7EQvO4ukTahnsffF5Kd/p3o02Z55
gaduHgCvLrn5uJFvsm6ztj7AbuJ83E5qyXjdAbd4Md4k3WMgauDnLZDqUa2s9ZYf
9DB38m3w35wMG2Khe0alwvSqCFti4tuE8KSjBsAQKiJaALa70Kj50l6ONtqCHXRi
IIOwv0r2vSuVUivMmmrohZiIHCuL2H3BO8m5EcgTi+oaC6XhbiOSXhmJccVNJtCH
KtAkH31ssyDPqs71REQF91cneB7FBI4S+PIStsL327TobJNUbJPYJG4h7EmhYIBV
1FCqmORyxmuDNxXPbeIOtMmKhaBcM+2+g+NAVedUiFAOAQeMT+BFGUPpy64X41HN
oBm8C0UTLlIPKCrewiZuN50/UUOGSWlRYDlOhx8v5WTF8J/bwi+pmvvVUoKnmchq
CaxCqXWmg56CH5e0Qj8qQiHd5jBORiqbIh75yUFmqQHcaMDCu0Vg2ojOz3n+JDlp
Fuutp6RQ+m7AqLNfQuDzDJHx0rJNb9jP2hNQUlCK17UxPYsqp2Q13qXMyDLtJ9V4
6ds3KK/oPnXECqHvOru1u6HJY+r8ub/0NgnW1VdVjzq0u/AuIpfXOM5m0EvxSjnO
fq8Ds/FZh9S4xG5tqXvJVkdWSJVYlWdnfv0eh1kEB/SPrhZUzOcEFMqQQ0bXe+M3
H8ku7HUEgYj++hc8EK4p8vmDaBDV6IXrMoGc3b3WGuVQCDSMVhdR+vU4E3X0O3dG
URTOk9HkSp0ipo338KiiwEq2xWStV6gDYB0nC6t+ThzYrYLZPmE4z9PY6kr6M+0q
UWlZqnZzA1Ahf7lSSiAoQZCwmeSqdVT5eVOtbzmMq0VN8+Pa/qoKopRtnNR8TBzA
/QWfQyABApra+GZaDRHEp5FGbmtsew4uyZCO7RIIIH7D35IyvX675oj0hCf6cfhB
vrzBcBCdIOeSeaHU/8bpEId3diNpvUL9tm5Q3Z1yzKK9qkK/StUzWylBRWLnI2Ou
hXKuvP43ukMXRz269SQ5kia+1yKcJwDh7mjtyfVjDs15WpPLo/iShW5tn8qb0CcS
qGru6SyWdZ/TAyj7+5AVLFZE3xYpn9DI0nLoB2kCqjakSx8vx4Na6BV4OqqxPumT
tfJF1dUXw3hBfS9t//DiMkXgK522exPPUDtksHwE/v4ScFAKROIxeQ/AuGSqnsvL
ksPFyVWMUaHFLDukBLf2C0z6zalSInlatjm2rQtRQLXv7+yzKtJjR5y00IMjFnNt
VbeFHDUPeQZq1ZYHK54yRT3kBvikibYeA8Y2EM26k33w1bgGfPzIei5gW4+qutDl
Cv7Wtc/4dkybtxigjxz4rGKGCLrSrVNiW6no92LXkp2Ia3M5Ewb52iEVSlKlrOnI
Meccpioq4KiNQpaMuBOax03ft4XHQEDLAh/Nf+PPFeNr481c4crdU9ZFX0ZctwW1
oSwMeewKO0iV/y90OxwJSNGVSCsJ8s7/WBb2mSmrLMwUlK3InedM8LgHAwp4Rhwh
D3X5+859rpYMf71LKrZiI2SgaJ/wT7hhvL1/nNH20IzejRPZVmwZ728F34ZjTmNu
lMzPhbNtziQRx8fkJtRT4nxtzHkwicsqv2IOwsHht5zVG9yPX8QvXnMUP2Cx2UmO
f4/GMK3Cx981TfIoSOPV75ZxFgI1ev+2M5NVgrbeOMkcpq6plaih/8YS8ii4Jw4/
p7mKV9F+dTFsIMXGXhY9QsD1qz10JkNapFUSRxrp19eGLxBp6jpkucksCrtroKwf
tDLU0+y5a5yT+lVjWdKd+dCO7e2ilkrh6Lplk5OwkpAVG9O+U+II7SC32hMj8oK5
Odkwh2rS35JoVTiz6Q0/nljYb0qYrLIaE7xAOCJVRl54FZ/zS1ir+9gYadZeN2UY
XAl0gYp9a9FMkNDzeeidg4Y9Mjto/5nRe8S7i9r+u6r9Lot6YgV7KFSgbYszCaMt
ZfZ9Ay5C/WcbpVInGNSCjaIXxCDbTs9WDzze6HcANNRzhAISgIrKmHw77PZ4hVfD
9v/T0Uql7x1lbGuLafriDRR++n/NcdWzH/kUqW2SX2uu0ushNuLQenW+yUtTjMcv
V6ebcTVxp5YnQEupAyvODopCrs6/kI66NX1a3PCpUhtUcyUnGofHI2gv20QmocdP
Hq7/0RRu4ua3Mo6XGFB5FSbTMTkT7z3agB3ejdlDE7kcIilM3Ci5GDNd+B0M/3lZ
hMhWI/b56208qz6oWSMlGWxwalJcADAHs0edQ6KJA/MzofqeGgtiCqj0JVHUMRq4
u7cnzgbgBpxf3dHupgn0IBwMq/eRvp0ck6LezPD+dxFMm4lPTfF/rlq1j1kbfGAx
wae+FMQGbeb1LXH17XRqwv7mK+XRbaD98qnZbLkY+64FPYKBD8UKYIMan2A+fSL+
LGCrFILYKuoaa+Kj53KYXROC84XkuCMA++xyAcr8lRs5mmoLrqzrCyAD9xqggPou
zfRZYPaGBb006rncLQ0BpTC46DK0B1UBKwTHYKgSwh0xU591a1iJkWKxmkpoiPio
9cAM0EPx7x/9uunsx2zLJu8eJy0ICrHihgtOP4dkkBuL9gnfRgvSTeckRLB6dLP+
Jk1oHbT0KUfFKR9F8K7T3C1e25r6knVan+e6qVKGY8ClCp7dm3y79UmaHiNd4+rR
mIVcaUbGpPUuRqCxzmFAg8J30s9UEC2CLWq4ESbKPaxm9dK7jCBzW6ZuOemjxgE2
GoxGmhJPGEqgxZg1VKjIvT2cVWFZMJKRN14r/3L+EF0Zv8BEBTBvDs/5FKkcMvOZ
NLaeG4DFUmTU/OzFUeSBYeQ0zOM4IvUWMOaaMsMqdqMe/WVF1rCTjxMCLRZzXLgD
KaIkGIwa30Y4CFsPt8u1ix0AkbKZw2AJ7kk9BO4xCQK6BrFQjPLqUHM+LUC2cBRM
t93XeZGTAvU9nxK6uHiEhg8uZo825QcsujKGNSkDhi2AjXK0b9f02LEs1zmEnKDn
a9tsZYs9Udop36B4sw7lISaO55GCOBhfJr5NDd/frK+nS4oL5N9G7RuJCd+nH9o1
basI/y0RPX32IUIrM7dqOcgsmH42/FzGm+KMNjGYktAkFItwfoCTfmJK16Tb9ngz
9g6aVjSWSdSxdDjvzQLuKrrSnp+Qoofx7scj9g5zxQgpau7eXplI5mTZOqyHQDEI
IQUM4Ns1fe+aHlIOc+ZtHeGH9npwigRp6ds6wv1BJqSCIFvPDwwNYvy+RkVwXz/v
/VZn8gekUcLFfsd5CDrxGa4NKIdUwNJL8eBX6x50rByP/yVmYWNLWeAINlNNnrlt
3+J/gecOqNy7MU2SuiuJbvt+bTyPbzkI1NiELDFwkceUioM0L7wgEBfdyaIJBrJj
cXt8wbcmM7DPhFBLMEufo2cV6U8IEfQ/Jtd0fPQz0r0/i50Q7Tc/VgIPKLoWf17z
ILBuhE4rrltvUJQKAbGniUUgbJGWQ3aZ+OFlUxMHcxrpBGeeZwA5gv4Z3SxZ4sF4
CrHPS7+7PydC3z/CyYkO3bpmRi6BMau3X2G8IrqH/THFi3RLBD9PEBEGBpIBX/xK
Ry9BQU6j22H0lhwTYmeGgJKvPpXjOpXFRw89gkQNXlQLs0sWBKJIRM937iO1IG3C
Avs47cCIDR9t+n10iqU/jJe+E3lYjPf6rj1j+UcYIWsdpB1Q4sFvTKqgT1zZknOh
0R6WTS+xOF8jsZDJNIxJgOtzL/fL5Dsf8IlorlPPdfxwPmbCX3+Ec9Rsm8Tgowak
UftTq72hiuncfzwMJYPdxBSWgkxSTkIrLAGYA2VYRZ6TEBXRVTctO/ahSiHg+UyX
gxMg4qpjWkwKPY8RVI3o3ELZ9BNO5S1y5twvusri+xOgd2sFzdZOzGei5E8fkQLv
RY8GzV4bIrLlmyppl/Zz3JFXLyw55aU8n8XLD6oCDxTHlOgEPWztC/+AmW4mDbAM
167fzmxymwe8+zpBgXSs24U4noQPhvN1WrtKwtbjBJnN5zuNqTTqfoXFYqD/0nnr
N7TCVh4vMpey0LxV3MT81q9rR7GcIxFeT3rMK9YqhhhiTTzzGKIyN57v1aoGd5NG
F/gEgsMY1D599zhRu363ynK7O2IL6w4hKtpCRVbTsQqq641i+XJkAocn5trX4ePP
plHKQlAYa64+i7Vr8rsUsRn4W9T3annFzPqUHpM8GGnEVRi6EKLdDeu4Mvo9zfrQ
VcmiIqc+Wjv5t0iEf3m+fHGvVLcjZhxIhMnLYs2ISeuYPLS+6uD17AVvCh6pWBLW
la6TvVZaEKv2zapo7dA/fl2CrceFshkBQnrSaRQwnoFmNzuFL0L28yNPdddKX38F
d7NWtGqX7VgGvEmYxVIOwI2RIHK0NUplXHW9rz4+uKV5xRsQzwk1+eHeZasccuye
xuq8kpD5yd69EXfXc0v9PbzAM0xjAgEIstpo+ta9lRdLP/1WP1QjgISAfvMXdaqO
6jXBIPLrtaHj3TvW6EgP4UE8gA78aoGWvX9yOrA5RU8mrqn/YmaD1qwwdYzvyza5
6tV9SbGiZsfhh7R5bHqr1TLo5z2wYfY8CavYdr7q6YT+fb2r93+Z43IrruhWqj7h
IckFzdMpQewyZj1udnW7lLjiuaVhBcMjpfyhWo7UoP0Cxl5YvLQ3n70x+le7emwW
M5/6vzIqDlV07ueJfEyqLT4k6OyTI4g+7PuAswlQd/9liOhVKoVVx8uHByRzPAt7
J5IbrdTTKzSHWt7gguhi3p0+rh/gIGBb5mQYyckq7P99jzxQ2XLlnPELBeTFE0p0
qDlZIAGEVH5j/Y2Geig5hU7hfMTEEjysDrXBq8FdoqQbC6VOvdxHNYYtdQvIwbho
zRhWStrfpuKi5pf2XArjigsIgkA1Rn828Wx1K3kzDJaQogrFFCjmH3nxlEW4rwVY
SsuQq3kPgwosZ38dkWFUS04eCecO+gl/SvIa8wK5Fi9vKAAKC7JuNizYa3xmIpuz
8Fe7+TRIkDc7NIvwWYQwhyKUgJD0IHCChvXsLtO0w1YZQpRrjkPKOleWtfggZAJX
J1iRWIYGLNeYd8doi1MLmZGHn90LtR4KHiWU0Kb0Ili0jxIX1rspPcjjzHkV4BMq
3WGknEv+aqE0ZBPuqcWiiXTTXTHNHdn2L8Tf/fv4BvJqrfNZ+4U20HfCJcMTYZth
0afveQJMjfCYSNaNTT+fEnt/D4BpA63eBDyi0LQ5K2Bi2fLv5sP+hyV+XFJC/Q1d
WZLbDVwCOEnxgjY0SPRWzL7J3tO53cRHwThfkyG/e/2J7Sh2dBYlnTy58g7ll4im
Z3aKs4QQESUR7fKaufKEuemXuRWKBzfcGNYHjKTGJonuBXzBcGtsrlyB9KXYNOhN
XPs+SNNadUeN9LBaULf+G5WOBxd+yC3cCk83Dk0ZRbwnWHMga34BHodgLxWvl4A/
QYGe86PJtn69khv2msruXZFc+1kFbUSGSjjhdxZMvgogKSe1/G8MYof4w6qpm+vj
hW4GLSBYinKiNBGI7E+0L8mI5ot4K3EmSdRuhcZG8RE6XiqXASSyucU1e3JsuOm4
fEts2f6F1AYmIM6zqD2qm2EfNuk8WSBJoeCgNY9I3n20V7lg2xvqA89OWE2brVE+
uJ84hnStCm3WH3tSpipAbSUM0JKPipQHdc5fTw8l7DO5gZwBubbQCvSyYuJVKxTa
qIaBoOMW/C3097alz2pNLn2cfWwgXxo9tc6ej/82IMj6p304b8Xj+qa38BJwNgS1
uzJk8883TU9/std1XUWJe4Y4fXg6r3tkRZVmqTkzMFICWqKrKoUm+xgI/5o8NX7T
WHzk6SXESUFxYUUkA9P4p8MSl4Vj5rPbCDLuxtw+wXIF3nJuBM8E7lkwRPiA1717
DwyBOQoKPNTjYok8Zxgag+irmrf9rLXvAiKfcl5K2U5aIWcniRkFwPslcKaKPIyN
alohtvHBm9uG2F0HuXC8XCjMeYfcxvhbnFnlP8sQ1ZO5uEv/REHUFoXBLu0Wh43+
Ni2hx1XN91JDeTwc3SNvhjDJVv95MMc+yIfJNVEdjEBbgsPvR5TnMjPn7hFHdvzs
QfaNbTFt3kwxZscgFjl4vPqSEU9btFDyNH/m3Dzk7H3RJO8r5COfxs5yFA6P0W/V
aI1vC+tf8myF3jMBGEpjqa8X99bJAFpyYXGdvmXp9XBpHdS/RIIM1ixxKMXRsZKz
79vqQ2xJpXEmUSVm+lYhNDTLTO+K3HkynP22yFOnpPIwsd8LqyGkiHE18cRUP4aJ
nHi+NBcqH3EFa5dBuL1FD0Gxzxl3pIsGxortSurwlCqsEn9cvuRLlimajsoeZO4A
pQ5z8ANiuIUJb8i1xJHjuhfXbimn/dttd+Tl4Oa8rUc47rUCQiP4E8S///mu+hjU
eNrjJJuJKpkwcBpNXNHRxTdCPrpREiQI8hNhRzcGdJK4Y1eP0zbCGT2H6EWynU66
PcdY0R72SBGZKRAaiYoZw8tzf907/rjr6n2jXUwS5RQ2vBhcVq/gsQGLKTh8U6Jk
zc2YgCC8jS3lwYjWYgndYx9rRgpFy+DvpwDKoFv96bRPn6DEImuxA8s2EC7F0xmp
+TlmDQc/Z/yjnOq0hfRpcp92VBGTNUvUWFAd/hLOUyXD+kuboqecsiiSp8DF1yyd
IoYib0QkQ8ZQlo8FYnzuOUSKO5BYuxDTL2oPDuYBzfQiPt5E6J8VvgxFW3Rjf3qR
yjjzpvZahV0r+hG3acCvkOBQUFHh6B2I0rp1bLpslNOLgiBTl0ODoX0/vNOg08TB
htVmKjNvKfIq1hqpvKECGzV+6aR4RIby3b7A9ryS9SoGVow5Ucnpr1xaq1mq5TCa
XPu16G3X7TpR+mMujozOYYGNKvPb66zgYqxGH9y+ggYALjae9krRd6P2k3tvv2K2
uGhTmSWY8JCRRbV4tc5LaUHjur3eZtxwyS8N/DnoRxGfwysbxVojzEanESv7UELo
iqtWI00AJaNWqvMrVZPtgqHNJ8v02i6M4EDxxTQv1deOloIpo/d2R293JnQ2Tbni
/nWFjBg/4CxOdDt15APacoWFhEyVXy5KPBzfrn/UdYBInm2OuzS741YowRyyF78O
8UyOoElcAZhRT2DFpcTDPCISDvSHqfSNUfH2jN2fSrDKwh2HufgFfuW/FrfRR+RH
n75QnohXmiXzbp3rzQ1JBP2uCm/YshNhVgTtFBOtgk+6ArAAVgHGU/ReQ3vWTtzH
zTqBliMsInztQBUF9KnNoO6qCM53T3ZIiXXViOmd9Hjyd09JRCt96/kkyH6MYDnm
XbNVseF70nXoIiellAajbZBWyfOBycwUXxMSEYGwYfe+iP7l93x05IK2rPCuN8v5
xotZfW061grLmiKvhHxFY5K2BdiFN5sC68SJLFatCXgqsi1vTc3zYNY+qJu/8GrT
brvVj1p4gg4cSJTt87HsXeTC59W8OTMKoG/4wZT9DSZ2GdAF5uvA6ycZDjGmUtty
coWL+xEEdVMVkkTE8B7gsR2Tdc/GrF/yUeCBVoY/i/efPjoOYlwqm8akV/qmMqWt
XaP09L3vsNZULjBs9H+E2DIpIihBe50cnBra5mlWWdzQ01qEDhkcoLH2sOTKUUwX
1mHlTR51BGn5T2oVQ+VhHgSil6L3AgmrfpNlWHLO8cbmjRV+RfH62LpQTamZ7SuN
mwQePLYOtNUWwDKoEo7SX+wrCKOs2ibTUwdPU6i7KAakdl//VQi1ZT2LwQxErLLQ
o+mqCnt/DDr7kHKUXo5QEf7ns2vSaZot+HVwMX8tYOOh0eHXJkPh7ybUPsRSaHXR
IoYRJTdGFhoTlXUkVyVDXHqHOzcVfYNy0wojWhEK4OJz6okSjPumvbb8j3xvW7oK
T0RbzRTGKU+rPUd9r/bkTm7UPTbQVzrKMbIC5LhXL7EsZ4Y9yxKeoY52vumSnFbh
z6mTXbnQHsKtGesurZcWYhs90luM2cs7yfk7M0RMhgU=
`pragma protect end_protected

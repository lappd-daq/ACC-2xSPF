// Copyright (C) 2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std
// ALTERA_TIMESTAMP:Thu Sep 13 06:36:44 PDT 2018
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
EIioEvjzK98KDNnVxjN4vB21lg1UI3Bv72wqcsbpeeNS5hxOcSqNNKW7+NOvjK63
0CgFPAozcTKU93Fnory+qNER1i1DnAN6tgkOyM9f/+BgwpBDx8fUxnjksVE1EnR1
/jGyI397/zM5neAKqRDl+rlFIPfXa126IcEX6G0IPRY=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 21904)
xz4P3Ly3I+6vYJ9PaiFS0s00+s27yu2Sr29BpXXgKHnp2h81OOMNXVo0z80w9W5+
IgZvUrHYhbcQrjxdYturcPi09s2zrkDCqjgIJh2rk6oU/NpDQjrPnd/Yl/VePe0G
/Q21TVE35jofEBeNNHJZOwPymLfyJ9ZdvUb7WkuQq0cAluMmdAgaCZRX/O2oIytX
7n4uAYL4xwxFePeIGY5NxXliq+S1RZKtCd8WL3fgb7HO3WFFXxNWIZrsY7sMawvR
GzfLgH5WZrvmswQGg+BztL8TsOoy8LGeSHK7+2+eDvEDTrhSzYe4plcr/SZVbAcb
c5+AJKLccDrcVgOQ6riao0RIr5LeYqBQgwYzo2ve74Epj4iMvCIeVhv6g61pJAvV
HJnYorrPL+iTKUHVviMnA00DZQc4MRtC/3TgkAWlVSacfE0bs6LS653pvs8ZrNA1
PmBKC6M3HQUkyY93KEZMH1j9v/HwemIwOaSe03dXBnfjKudcSNTKFVzL5M3ID+Vw
oJctM1/onPcjhWPR0QbOGlv0St3nfJRIMCdHMZjURJw5bmphs1Jv4UDK99qnL8nt
TopWTua12gUrh3pX64vQEjCjPUxHzFSlVwL4sZtbexgV3HIaLszE8Spf0r/Uziip
/lVRzuRWUyKbIRqpUNozaj3m20kGU8NLC3Rc0hdX+KFoSSi1SUXd+jRZgwTA2YsC
tJst1nzZq/dQ7oJB1M6ymulf6SwhpFVDjA448XTcva8o5tIEY0taaTinEiIQVlyA
1iLC7wq4dts4Xv5qPY9oj95kvt798D6Q2G6NQtwY0a0bk+LtaVEjO83oW00Fv/F/
2yAG1v1FHk+ti6QLIDogYwqbSG3vAMv9sa+YbqCNeKSGgd7OmlotV/lc1Ztu8LEy
ene8RjmSsb7ZSy8o8nkiRDRx2qVbTESIIA+kk9adkd6B6TvHodrUtWNNzYb3yIc6
mVQpbxLVFnQ7Oj7d2rWQEkwJsknVXBysJ0eQr0+OpwuxHFsPjsGz68z15TQzySeH
HBOcTZGhiiTI/LisveDOQwj6/CUiaCjm75mJft7DJ6c0K/3DyB4dK3kd2i/jvhmB
QKa9G3Hz3HSe30izgw410dsCBGu9DANCEL77qwueOQSPhTn+YKIiTxJMbmcVXj+u
KUUy+HlY1hQ3seAm+gDZxE0cSmaVZYc7Oovesy60LotOl5T7zesJ58rx1nhynbg+
VtjBLMrwv8rtJFZAsuIVcgyXim4w68KqKDY2eX7DNg2vNopwTirOGVuOiy9HrHPA
gk74+2Ybusq8eINbWzU8ylI/LOxzAVvW3HBz8a4bkd/fRHi5+9L6mMLxFVoNUd/k
BsQ3V/NrzHEqsliBlhgoOJf0Z1Wir42xO/FnGPkkh5dcgCPV5pBnxOoSrAynENTl
+6iJylkIEZK5D6pe94/BZLyhvco0Pk20L2RfrHU8dWu8SnNdX1Jph+8tJna0NlAG
Wtfc9CLNH3KrWi7LCp8BdSMKRSIJnGiTTtu5pw42XM/JrE7taZZ77pnnGyL2840K
sEsuKJ7VaayJ6WY7Yf9RCl9bZMYvH7Cohq9Qt6H+GGScoO4VOhf6Mhuo4OyAnXM5
VYbtosOqyAbdPPEiS757xfoXFeinhS0pcOuv4T2/ZSAZdCpJSbRHRCV6C3GWeufz
wERGW4mHq0wc6pB4DbnfYGVCiOdc5R/z/vJVhhZ1J/C47fbJj5q8yxjko1p9mIeZ
eBiUIjupkxJdg1/05dMPrTVMPmoeCwaQ/DBwneWML+Nu+SSQ9T8gReOMo3vqp3/2
5MQVsODliTReI1sm/8ThrNNYmhbXNxCg7Rw70E8GT4ILsvVQ2mTGnNsqTwspiK6n
wZA1gGrnwQEm73CdqiiiycYnt9cnrplZ5WOA8kUa4j8FxCucr0xhcXP5blTxGwsX
xo96HqOU2j4yCiR21acfsk6je9wI5rImrVOgLtzDwIpa1Lw6XkJNiI6kztqw9xcS
ag4eOexUzZHhI8YbNWSPTwzhLguVvsVWS+4yzMizeagPQsdTDxLmaUO8ZNLAKq5b
vOY7rbBFUMcG4I9aog01cMcxSLAVgLhfUJ6Rt4N1sAJdELwWMtKdbpBJPogFQqfa
+x3SimX+z/Ak5sSx3ClrKf8dc/A7uRcYWUeJ3JCIpHKwVCYs1/ZX9mRAk9molFLf
oWvMgtyDHBDDc3ZNaFxILj/suq8egr+0Y5hhaM31hvmUEWYSSV6Z+RdczW06t9KY
BaQg7kUljTbfPJJeea6Xp+VKsDAiUL1N/IEQlXRO4tFAP9AkqrF3IXWIJMHRjH6W
eK+8plwnmlHicMnUnWqA8vSQ8/0eqKNgZKr3Qzvp5b0Sss42XisbQS23R3e9+46J
iA4c0hSw6EYvjBwpN+R3ROmSHlhYVSsEgg0rr0n9lOJNF5UL/BMgLyT3QFVY3rUc
iQsh/HzCXNCfandQggxKeAqPpVX6y6GCZ68WgEdQsv5eoajM5JANWvL24KqQEaPm
8uLoQjcd+Atei0ikADLQRWAaDOeHOh+Qlf14HVULHKU9misqwoTqbIT8XvndttLC
RmbgDgwwjcsLxysmFmysXXWUEX6A68tgii+C/9Gqbyd2YnMmwIr97HG3rmDmDb/y
7YosvF3eQsp7U/NIdpNVzPo+uRN6wq6Eo3zNY+kcj4gpdSbzFMSquICnNRo9HdNy
ofUi9VBxwcNo6krX4KufU7M0EGqzOD2zfd6Zjd7a+7yV1XtqQCpKY7kPtbNdeUZ5
Bf8/s7onSHMG7SPAXJ9GcZzhaJFKt8Wsh4CEFtJNatlFKeNCcd0UMWxZPWpGLq32
5OhKJAVqC7f2eD3eJhcByKw66ufDhV5OXKmsVuhyR4Dz3UQ/YHNE8fIRcxMP4Zhw
YP0zG91mvCqe13xd6OHu20ggFDkKMh6pHU1DeyhLRlGqjfRmUzuAm3pcNeJil0IU
O/QOEiTNViR4X4uCzdr08/5yei+nCP2k+lD7GvkW5Aqmx8rRN2fyNg91aDZqZhX4
j5cwA2hp+03WauyL0CVpTA2Tws62iz5aiY4nqZi8mZ6pfO9fspIE1RRbLQ5JR7F2
8/8Iykp8zfXdJDjKQczDVCnIvH3izZ2WXJF8EJHvCVxI6T6jTUj4l9t3RiyCamMt
Sl1ldX0b8FJ8obzL4pTybnNBjgqjKwrDHwofbMem80jvbmtw7AHEXcqMI8teGE+p
lWIqCMG67/MeO2JzO/9h0L0iC8mjaTh4W2/USgkECzPxDK5BCXMxM91g46lmw5U5
w2Dd3GyBnShLJbnx+Tul4WfY28US8+JW3rGMVpEL+Bwsd20UnjG8LiJvTcb9qRJ9
SL5qV7FRMb6BipvF3HHCMnbl/AImVFu/NipIXI5S5n9fDzDbioO3rwuHnL4LxFaK
imYI/M2fJN8FdQQmB72Z4/C17KPNbHtN9jIPkMEknHYMM1+s8h9NAMviVhaIvYkq
gJK2+c/4TYREECWKsl/IH4dF5a6/3IEl4j+8VkFmeAkqywqrGeOi5lj9Xj8gIDgf
RKWV8CjVpV9HGnBVn5lRCzTwT6O2GMuHcAiK4igBbx+pubzCVaQfZDBKFUiLIkoO
biXKbLiFXqPzYw4Cwo8tLXas0h6nU015DXc5qO4zYyq1NVfKlMhD5CYH8xcBNeDH
Gp1BpDF3Cwp3VSY/yca7ApemLz/IltHfO2KQcHmVJhMQHCWSgVwQ2mRLG5mtYEa8
9CpytVbAamFihowm9kWl3vmX0Lek+sJwS871txXBEoL+eWaKfI3Wl01Dbe51eLqF
cHkiRGJ9VZFzByXC5MXjpuOeBi57cFKbFNwrkJO4GehWr+7ZKtGmNmJ/egy6m/nL
0uRTdKlqfzdk5uFKFa7rIPVsCGmbPzdHVxq7iIJmnZPyFTxo44HkX7Kn6swA89fW
K1Dgo8WmbNAQ5uNSitqKuA+vgvBhbKjEg4Dk0q+0Md3dtv/mjspQUxz7ti+i0jXV
p0UN2uw4ze+Wt29Sa0wlY6Thn9OYuo4Ppznmsxl8tvUOHhaZxPXo//M8sj7q2rBI
CcbWiX4YzK5bshLY6VIEDaVEEGp7rVtw5n+GEn2/lwv6K9d35LAw+bm84zPx3Cwe
WTgJ1tWHafO6A8aJ6k+xJe5n2FWSb1x62JQgcfG4jMDZZQ3EeGi+KtLf5tBlia6l
nQy0c+4uPkX8A43wBlRwZxXuO1o523MyenNmNXgguTv4emy7xlyYkIGi1t2nNWL7
TCe8dImq263qG2vpVtiv+lIZ4G8yT6adX9JhTuA59bz13p8/Fo8R9rKOsLdQ51AW
50c6cZ15r4ZO8+jN579I+dZPOyA10iz+UhiW3hKCG7CKcRXq0OfI1ag5X1YlMwKx
LYZSpoUKT0XjgcqmdtTra/FSTjUzf57FxpizeHzjNPX0f7Mk0wG9sFhrporzE8UR
4UorY2YMCoGfXHUaMmhsPOsE6VbKgY8vprYCl8krSu+dyPRYuqgVTRt2ic9cxqNc
taKo7Zhw4HNfbj6pO0zy/2bE45DkPtnpt51Y0oZB55Q7J9J6P8ZOMBndh9oXcOx5
JfeNMCEszDvaFaEDdnHkucDzXd+1WU+RH8lvkbRKLY92s2Q6xji3lws7flTLRjBN
TrTdrgBOJmKJZmiToUNASEtVepwGvzS4xnvsiYbP1iyXuFxQpqE1xvhZstC+OShP
TueALEV0Qs8QbOP9VwPi2TUngdlHvwH6/1TGDz5qJq3uwnVRfWBbww6EWHKY/XFP
cfHeOIGSr3SBX63eQSCiyCqUDYWLZo4Q0AjYMCVSwJakoDGkLZVZXnOy5vQPbzbj
h2pjcXJCxLeZI64rIvSyLn3WKzJ3jeVNZolX8jaMcjU5sDK0GuapUTMBpDL3OyrR
rh8uzpB0FoGD7ZQnhgmuoxECrZoMh4/jPx/NKume6l1QNgu95WBgsBnYyveDl9Ws
wVO+s/6q8/ToBAQmhmGp0zklhOFyHE7DAAw0Xn7f2FOgcxvJMH7/g/TmzXe8eL1V
jkx75E7rS4FzliEXUKS4EgOiNKk1+GO6VSCu92PbvwZ20uj7NluWZ6Vidfdd4WmP
zfGWwQ0687v0pL+KqjDGrTn9R6/0DGmbQn61suusqhNZ0nWLlSxye+BmZ5zakRPC
dyoIVHy0JMYRlZ7xgiA4HgMg2WLuGZraGLdWCgAho6saj/H9+pbby1mMGLWz5Qor
b51d1iKfWMrkEUchSRjAJuUXfJD5kjH4O/ZNtKcvhf7wvmTIzXMiwsccwMLVOTD8
djJmiWvZRwLBy4Fs3Bj4vr8m9E9OWol5x99xKsmF3AGUrmlh+3Hb3PCuQBRjtHvj
r/X1eUNN1oQOLbDTltqGFkJfgSjVKGQbWpcYYocZ9zkKdQ04LBN6YmaWDl855kIJ
/uDexJNujQixjNpN3YYR2XfwO0rsulML9YWsfrXn6zxU0euwWp7djasfZ1yD4yhv
tToxI/1NEkqGDGSobWJMhiV/rXyr3yVRc/hfrkjXmLWzZFHC4W56vUeTW0Ds5S6U
mcqOurcjCRHCfqyxtMCdtvwZkpu+p/hJ/dPrd/WiVK/lSas8Xu/VTd/EyBRDE6WU
/xVQEv0/NP7Hoj+P1h88rfes0yVcRBGLe9Cq8f7CP3YwUdjN6Z1JjHdUhoapwPjM
0ujT3utM6PC9YkmIU/84UHX2XhrXCi6gHlEYhNRUQB0AynPa4OMETOLfVHxx6DKS
MQ0q9rSLxJJEUjlZTpD6+xF1RJe8raZ5XUcxZPmyQq+EmayxI+h3E2WZCbCATGhI
A61vaksD9DFJ21RKdBh3AOwkvVx3wZrLLQ9jTwz4FALV1zHUVR+y64KDJU13+BxR
zyVCQfKGSvtEtCCJnLqYQzync39PHOymO1EvlpcXzFmg2jX4weJzSEvL+D3t2mR3
ps6wONC23SMI95asYNqnzPhmtcaj+Qckb9NRj55NZ04yJe3m6mSGXC+ucdThIyq5
5Zqc6HLEWy6tzSG5BVBBnSYxLjbVjqS7lqZFD1pKUObKZH7SOuFSy4GfsyboxJV+
V8KmmIP9HfUShoWBv0h3fzzDW6/Kr9mRTJ2VIfgIzdYWfodmeaVja0Joo3bEo/zg
NSc12knaYUfFe94HH+ZANxxpKc2YTfs3U53GbhWmxhnrVZ7d0yOuYR7scVU1vEtJ
Ot6EH62ML6xPazXY4YHymPzfuUagHCXIqFLmi212D5YHfmAYcn1TSxg1EWriq1QK
Z17QfUiJXKp4blGGiGBjWSsWFtLUcaRI2JCBYRKIIQCZFboP5Gsb0cZsYMpmdVOo
p0E7iViiFP/qpHAfzXItv2CGmVsPpsGQnfLQ7wGZ1tMkCqGyFm1ep9hWctPbmQdk
1+4Zv3PSDYIck6pzBFslTCKSWqL9ToGjvfk3odtOWYWWBXQ+RJbAYBVPw8B3SC1t
tyXOd9Fbvdr1wRvA9+MUqZU0OD2Sa8yl9kmBuctdlyGxe3VV/1UI0xU08EOOoms4
ZhEOnw4PhuhLX3ZwpGMZhriK2h/XEOJlu6H2984ys5mcYFI7zCbGvByw9xwr19KA
DnxTMSkNqMnFdKo3Jpt2zG/ek1uSvtDNEVCdqyt9ZRVOVT0rDnWgewv5vzl22lr7
UEwjTtU9pArfldYIJ6cIOeRvQ5DoRS3RJ3xEbGMaVvZjFiKaT+eRYfhiKxNsfEPn
cCddN+1RTirq2CCSBnPWYnyxoOsMv9nFa8hGdDR8hb5O2LJ37A8lvPG+CoQ2co8p
SeQxJ3pDYDhGi0QXvnYRzJkH8NlyVUSmBKDftM21zVjnhs5hKRArKKgrYiBvUYZY
/prZMli76f0YxKz+tDHHIQLlbzpe2PeT731EOYgfYgONgvYvs3Snofbtd0NBBXUd
EqIXKOAqmiJgDfl3F4MiCUAXVVtfoLvEMWZxWzkrmLbkLgPRVAjn0XQi/PZqQQnj
389R63GHwD8ThxNUW2U4k5tYv+Bubnv4fbr76oUURTmeL8r557CoUdAoaoVsKdBP
jHqCo2I4GHjCrL32HWwBHReKfG46UdTqGx0YHsE2BokHKRDV3F6Cng2gbd+ny1zd
TTN8DR4Sq2MmNCZSCL4syYrHJK9k3SmFybnZogzkCYGRVV99bPZ1d7bYxXAb5kRm
BnqtAp/IgjP1Qp2ei0B+FduoQGRgZX3kajA9HMoTLkelWOhQuAOWdx1DLu8k16AG
lMJqojwiJE34BmF5GeuhYZIR6OFOld+ERohUNo+Wi9mogbIEunMXBspjznRXx0Fc
W4KnpOM/W2n6V6RZXaug+kwqZpWkYwmvaq3jayqLxKFSLm3b+gRDW1xa1BzvEIxl
6Tsn0WXuse/QHEqeZSX/GQMFLWJQBlFYyYQgDhBWYsJ8zd9qqaQqdslX6zk9S+sF
63IgOX6G8U8XPbSwGsrqsv7N/Y0kNBjHrsXsPEOkYxXANkBaHkzs3tpGxgaoG0of
5GlPCMG72kNfyKx7rXU+18Vzxb3FlxLfeXvStYZdL80+uSKrWmqCDjImxbgHqqGX
riEAy0LaCc0fiLGKDU0HV7/tolvY8stOkjMcufzS7+VMx/SqoMovxk9nKRBUxeWm
h4mo2AmtKe64CFyeGK+ncQamR/8uiVfIxmNPYIc1ikI9FG9KNS1zVhBgaKjNz5pv
ymT8HJqFUylwprZ87BnusY1hLqnPd1tXQWDQX3luPFfGiL7u3vBAIHnK6T6kMyqV
pInXksrF+1gQPB8IgRCclJw3RXrl70aeJOl5YR3hlIG2Owg/dtPrv7EndSrlKwzk
s/3mwyN8ANCMB6Vij+XoHot/ZfaZWmvn4M28ZHoNci6xsxaVFeq8H9CT6lp0n3AM
LZCce4oN56meHusfJOH+dPem+V3pILMoHkAX6+kLRVxhc/1W1pjpEXRTacs3yDBv
+CXXoYLouKlQr95Irpx+CBr3E8fWr6gVaHax+VdWh/q2oaUin6eY+iYdSoKMR8vJ
QwHty9l6dE4CmzVw/9bX3LpyYJsH32gEYcOeZwt7RMWCFVbTeRChdGgZaZ045adr
Ww8pxJvNZ24wRNp78720MMjSogz0/qA9jiXUWgwAt2onvKzJ9swUpgYHZgTcK480
ZECUvzuf/L8Z/I+pbqpQSeRZSQlRRjLn6zANLcyPnXDA4Hx3E7rabpNcQNwKHMmI
P5xBm2XfjQHzfdmHEDQnLC0AAfxRagT1dLxf3LvWS8LtpWJx1fqfmxgaqBhbu1yF
B7PAXzSvwKnRTFPH2VE1Ds/CXYbjuWKvOa1x6cN1dn3bvS87MgUPuvJff3lVVAxb
rVSiE/Yan0I/1585eiAX4ts+MwHog3Z0iH/6gqwm6KlZMW9sez/yk4wimWpOu0AM
X+s0HtTLcjKmPJOQq4xumbi4vxdZ0p9eDHFcQZ81tkujgi4maOBf9AxlKgFRPtWx
OttqD/5yfWTqGPrtwFphgK5SSJQzJg0hpz+gUSq3PTV9Hbhu1RHy1MjxYZEAwJcI
fo5o3u2wWPPwcJF7vDX9AC4LPJMI6GRSsX0BowgPFk/1LO9seY5D+foSNsIrn6U5
3oHvJZ5uD6PqJxHD2fIV4XWGgGZM05cu85NFFdTzCE6VRTMwSQ+fAHvSLavROaGc
Eedu3PI6itJwkaWY7RwnSFsgNmJnDYsnMLmzBtpiz+i+xhS2O3TrtePnfK5gxjxb
mV/iw793H6k4AUJu+oaP9dabLcTv0lVxjeOZ2ZwY4NrELK05vZ9QlKkx0tojDD3f
gU2a40A6TxtR6wyj+u+dlEQZg6nMTPz2aE2y/tyJPB/ExyGwITomKhLBX/dv2m1Q
UrCL8HKORf/4h+k7IXxrkuBre6r5tP2x/KW5sXaEo9uZl298BrHziUo05VltoNKg
UM06oom0tVPFAfZ5YhmUrBxvGkc0V308Ru0GW/VFoUOHlRBjwu27RtUV/0BIHdpa
Uo8CR+l0z9xbD2AQzUxa1mfoDzJRE4ntFzzzaKpjeAAgaY6JcDDBqWzpd6M8bloE
e1Ab60T0I57Faew8Byjkr9yAAIzN/YYuPCFupWiS5uSv3P+Ap3Cgg4+yc8Y0+/SB
6ixRimEYzsh6Xo94q2D0PUyluSrWO4mXKkNPhxIu/SBeRoIlQ2Tbihp8ts4yuBWa
hCdjmhAq/+9cezDU+1/e327W6XTc97s700zP4oc+n1G8/undZpkMifp5yK69RZ1Z
9jCLYrQo1PQIz+UAAd4LU2UmhYrXrWU1ztd13qtxp02ywAL7m3TxuqSOa+/iY//3
UHCqccTmvWizUTE4WAnMfVEu5wbFWJj0msfXc+yNId6GdH8pUr/ZNKL/s6KVV3v4
ly2PH5uRtKLTvPU4AvqmBszlpRNuWwwD0D3tYQ6R7mHhYsjFnSNtHtgo69FeVPx0
q3ypelzWvqG0OtzIxf2av1UjZ/fXzO0oIc1NN1vjdYUb2dkiaVm7zrcfm3sztKB2
Qclru7svCcQ9wuKNV2A9Vwci5JYE9JH7Z4wSpqUa56vQWAUUeJqRrBB+UwVJxBVN
ZYNHxts+3EgVJk5XOiXo4Fc+qxtA03/cfC0eq7F5duWf/UOulCqsDlM6Lxs4srKN
b5Y/DF3ltwm09H30NGFSm2WID6mmdPd7aqhEQfLwzLOAWHlmgsvndyoMEr0i+9W8
Udmfxsl48h1T1ieNzY1qPQcUhzRLR77EBlfF4mnPj6lweTg6yl73eowypwUiLRKP
QnSPnYLwAtkSyMuH7nhYZ6V0juVv262g1QT0SKgVd73O4lGVA+o4BN9J0d2EUexO
ZkspgrdMa2lGJK6Dl0/7vbfZzGM8VC4HEKUHpSSoOGx/5ZDxE+elRKlsa4Hc3wcQ
5rlMO3wR8r31BWfTU1ZSr1SDB8UAJ0CY/KRFSEEUSptN3Ei/PjH3s/0aCodlk/ux
woklgM7Xz4VAcD2mxHuOQlE3zumA8/BjCNwnOu4b1Ni11TJyS/k/0RzakbGW+54a
G11Qp1UG3Aoc3d5S0APnc8ucQHqbfiwzGyzhUZDs1/Xiu2j3QwCzUpFoYeRf+IhJ
d4c06ObGVrUpV1nNodMzfO51vep+dvEdx38HPXEJNLaKjS1ls0r46FpNr+h+gYaU
zcXQcOJwpP34G+yNVqnuYAMI/hwtZSruNBt55CF9SpvIksHSR1PmX3gMpYqjJueP
2BOKaDUpTbVLD/t7+tv4CqxJHK5XM/MHkEWj71LAjzvcmuD51R0WMuPSli5JYv3r
GRLBiGqIr/gtKm5Cvvuger3sNDXAkF+yv78vTFYaEx+q/eMsjgHH5y5gHcbns0L0
U6nOBScUItL+TwXQBQ0FY1SZBp9a7Kj1EBPcUgKHjMh+8x16TvosRNDe4xYw4Tn7
J8xpMiyL/vQ9g6biIX+AdXSSYL1PYUDQ2rtH/qQUULnL8cQnNcSQ0/gklQRvBthd
xyFR3hP6036e4I/kDuw+WwT/pNxMSnHwez8lEBzQwJNsjAlAI/VJPri0A5h+hxVT
aC4jqCrwjnnQclskB6ccl84g1Hms0czSTgeevq33m+TPTxlReAoi99Yq2jdQQj9S
2cT6qUzwn2vUxW7LmVafXneJCVAZHmcKqglxX5b2k+c+yGGKB3bpWLlnH9w6nJKO
/HwE21IjSY7vVH/R2a0JObh/tVPGMoWelEEuMCtQTg6HffdoQbP8QeFy6Y11J0sn
U8NwdWP7dsEW0Ev/Zl3Nco0uzVmlfW4SPwYOsjnrjkIjF+A2VC+4Ih/+rjYe8qbJ
ExQSHGGG8C7pFnIJtlAIew9HkmZBkGjAxg8Dz5OaAwT4ecCwx5tAw29KnDkuuPnN
ZIak2TjDKM4a5eB0xN5FxmVX4MU8KriTzqy4BK+rTcI4/eHP5ludfHlHH+cD9Uk3
U1pKvOAonE1K20A15XbM6rtShsT34HnMsUvUN9MajZSEIUGRfjfeLj60IvyKWc/a
PUG0GRAlD0sxCl1o+0Z1MqVb5asHqB4VLiWHLICbFmsSbK0uK3oQ2Jn67bjz5z3U
LwY6hTpwBVyoyoNYUgTU+b6wsi8xpp1X1+f7VmoyGuCxT1O0NtAarxlT7SIJ5BXj
uHsFZPIrE0x3W0IodwdzD3UjiyIa3rCmVstdt36UJFgh1gmkirsTNJ9fH1NkqCL1
L5JY72Fzb3bAZl1TpvzdjtLoZLH5bOp1CAvpEUbcSuGbRQtz9QfxgwmxG8mjBeTu
xw3M9y/+4eLPP/1DWtin70SNFNK4C7FvdCVb7nUGYqzLIJlE98vcZkqiEvvLdXEM
VuFfwDDxeqr7pdcawkPuciff494OUHz0Ojng64InsKHclV3jOxtGUy17vEnVwqd8
ofoGLqomFaqW2daHMr5k90NV569nFlLHjWX6mnLbwOwV09CjcIV1xHSB4s6Ro3/w
ZHzXC1JtCaPh0R5fg9mY5NXLEQcSGy4cBiSkun7crSdix8Q6MH+XnNwXLYD9ec/h
EsLvfH1rHzXocQIkvom1o+xkyrm4OKgbyOB68QlR1N9w6MP6i7UnGXDjbF0P/ssv
trO8w+BQdZXDayGb5wEVUNNdPuVTfqzNHBjm+Z+6KDUHHGIG0uQtozIv45OTyqAr
WBF8tQGeSEoRUio/jCr1vF706bEoaw0dzuYbP7s92qCHL5jSHxiY80R1N8rcRJ5M
14pmci3NiS/eexxMvMEHgXmIk6BmMoOnDikmA/yCZxFVB2G4G/zVLX53R61xUlck
qMiAgKJeC7T2xNiAFjMDNibeUjven6CLNxgETUZPHqlog+OwUZDcC4UPLEedwuXZ
U4EJpNQc8YARsD9I+YGb3T7CJtcITYcRuuceqcc69P8p/thWOd6sUUCa9XtDmy7B
osRWhjM/cR/VRYjJ4TcAak8buFJdIkV5wdCP1/j1wDsG9dnX7BzT3Rrs31M35SJL
DZl9MVfhusz9k/FZrUAwxzRZGPydoA0npuqwfl+Bv1PoE3LInXgqLFt6pV49l0T7
E0VpdScSgPyNz7ULuWym9yuEZy73Qq9pkpNutb1C9+NU9+kufQXO3xFxBxIvUb93
tQMyOgqMXU+m5dvRed4I/OzBAwFIp3yDOFMiy7tAR9/Zk6WNOJT0IiEzKrFM8Tma
JVOIeclb3Fzf3L2UUuWWkgNw8hiLYnYoALYy2P0MU0XSW7XkCrEdpXVjD2oKU2f8
wHawcG3FV7euxfOWT4PQrbtgP0VxsTsvRpDHFDR8TTNHxHmpf0zOuO0UuWye0aWg
yKsffHtJJsiDlhNRuMODlivWJ4hBSmU7Gki4YtOzplF+Gj+J4JHmhsSCnfEIMIyf
56803gUGUYyiA9JanoxRjnWe7dIF71lt5wBtc/EsVPhqm/qmJ0+qZ4fnHRUbnkiH
iypF8jglPNQ3PNvXo2s6Ws2hoviGRxOVgdaeOhlx8wm4SkvHu8XYvlDQo5QAw49a
7OBT/8S7LjKeYm+iLxSQfyJ36sdb1CFvWE/oE2M1iQzJjWlrpg6kkDCC0oS95lMk
gRbiAMJzOO3hwt+T+mGMzUiyzyT+NnbLsR9lA8WxokDBIDIeQCeMrMj7AdjM8Ht5
OB5sNFesZkeeiXJ1+TZGe2OBRzA/k9FgcqnsvDG2QoCCGebG1v9TXBn/EdE0cWDN
i/wMm2EwQyQWsYG9Hxt5j5UDJsCDgFJs3j3AugAIKVmUoc8jyBk8IGiLjHf0RXHf
R3RapwLvB7vDXZJQ+bAd5nazWItSrKmq+aj8kzPpOhYUA5PlX2CnV/qeK4ccOw+u
Ewg8IFSY4rQ6q4WpJqhs4keOKpOVl0XitnuM8jF+Two1hY0t5eHceqOjRb9YEVBY
ZARi+GktM0JZnYBI0j+h8lRO0ocXa4fVaa718iIB2fHoHlrI54uqs+4Jobapl/yB
n03nJKkyu8sU3l0BpG0HR3sJSp4laWCv/SSiSpurZTlldCfgtSsbfflK/23wYO6K
3VocHhEaXdV0xNSSU+eN5GLubTITr6KcEQpGoqkPrAmf7zDrpAX1DyEYL4ZedonC
rrSNGoj7NoX7zCtPc5id0QGIgEUu5CdMKM8hYF5LdaiVhuhyGZqbrdWHC5NAjQhW
VVoo94IXH2r25xOxIT7SIWukB4nQ8Xlp2FkgQ+iZF4/fLD1h0cbAQ5RKcZWGVurR
sjB91cdTro9GJFeq32m3tUWVTT9epxDXQRidXJ8NCPZiNxUt4/8IHWKwEco0qFT/
YOe+AqUOBrT4pBYEZ3kjdHk9f54YjkRoqxZef8Is5fW9ffcNbaBQEcjzksQIh2Jw
FCQbXEl2s1tuByq9v6M+9wLCatrpoWC0e00UR2iFMNcLgwgA/oB/ebU0gAqIuNEo
vKNiki9mFlPBx4TKvKScaIWGvVN5/l9JBeXIJ7STSQwY41CUa5JDzFTlUxWA+kmL
gJM/FjgAM45tAcqZnJ09x5/f5AnqCIr3XO8kCQdj2k/AXJ9AV5zv7FeXn55ge2oY
loixQylQtY2VjHRpY1N0cUK35pbq/w2DCQjafMCFNfxyFOPmCAORhIHTzvkgBzsQ
+xaq5gy3ualJzrChMEJokI0Z6fkxJGaDvBXoi3HDFVFWv72jYRSl0bcxnk2jQ9yH
K0xFLG5m8NMxUUiFYqT4WPVgijBPi8c6EfZhiD8xDE/ZXKds1JEiQCNUV6GyDXz1
rkkyrNOv/AZAI0FkPejWfyPOZytwRggeOnZwJ8FGRs+XecgRIrk6o7y6KnEgZhuN
To+d6OZX7KlBqAO1/2nl04IogPM1evmsJgC75erMW8nmkVC8QMiDusP7ilzhQl/F
NOB+/BqyDeIy+Za6UkphQd4w+BXZH12bQCRsLaIG188xhbPaWez9ofcnyTW9vR9Q
1XJByJUOozrWXjOfF+q4gjA0ZK6TfIZf4H11Ak2atePvgjsg6eiA5Kbn5OlJKN0t
V9XgJ/GelmolLG3Fx5QIgzEJq2Y053KJlVUX77KkeMC6UrDRndwbz53HPhs8IChh
49yDRxr17LhHot2vegI3ui38TQweXCU64aYOn9Q8eF+LkCqxs3+GMNpi0pjkG5rH
WtGdKwAHbRB8qBOslaPt+OFSe/FwNly7SsMvrA7XaKOxk3bQnaW0CEJ/MpJFyJQ8
Yy1O4WuQ333wD5v9C+UacdyKMaxUBj6bxGhd1zpts7xmRy+ioE/3raEFAKcBI7C9
rpMX8VULP+I8pBH/bKyEtpXPHmVnjns8/bWLM7E9aAq+MehThTbJCkpuIJjuOK1s
lKyS9RBsVZUponV/1jffCuDlbvIpLsHf8Dn6KE5WoC/NoXqpAUgeRQuKoIaSmp4a
oLMNc5LAOcnJ2NPZrAZg/yTVRqxFhNckUJ+2JstlakZp5lSX6rdtScP9RM6q8LIs
+oWMgbJgebEujeaYCacIk3dqmoYWbIT/+/E8fqxjNWD0juZLnx5N/XoilpE1mo+4
ywcjyUsYKzITzvFVbpvZy5kErTrsJBVY907846hYRJkCvc7snQObDxZJIo11gGP6
KxHzwHH7voNSoIKytEWpkWMUwYcwJrqhcuQz6JpEWxA+Xi6aVQqWVjRXWtQmJsr4
cuNYPH6QAhvLaY5OUm/N60ZKCHtTWhurnhrIcodMdoVmVMFKJceo9xUoEgnGtDi/
ESP3oMsRWJnaFDlktV9iPGcVUQIeHKgXqnqeWa7uuBKwAtHa5g1h+vDgf/W5bmRM
MYS2SvAtqAhuDhskH4cDyKPTmp3xSB+5+HB+Ah9vHSaGW6tkqCwz58BA4kBh4kO4
/vxB1kqM7xrJN0GpeKlPEep7U1+HU7sGU6TIDlWZlNpIGzecRDW5JHC0TIYBvTZ0
jZs4FKI2fUV4a34TtjE0vySrNmejyj8/D9i8U1BH7NdcDpLqC+xNpXmMwoKVfo4q
KjlFieTYv3R1SWH61eB9OXrCc/dfqrD+QRwhdi1GQidYuojH+9DshqoHGDaM7Z0Z
uHg+P9vY7lI+YtF9AQF20+0cEz/So2PhWRcxPkNFRdQYzV3Car3OudYb7uHH1H1I
8ju5s5gsUH/2V/RD1huq9BqPF/ybpreA8WWu4VlCX2SRCHWwBjAP+wbJB32N0qOt
XmXSK6u+02zsR/n5JLzFnM1jAQgX2LA+D5IsCf50YwfMZWB/aUppIQQAL0W9JJ1T
f4FrPJyZo9Tjq8IrljQhDbkeuuvfwSLs/Og6zMP6fR1L4O7yH38SdVsgasXoBbiy
/cEk6aMeNVGtWYdWo4OhroC9aV0JI4VHP8EPU7YpIeqDzwbsi9p1kDs0swot7IIA
w/gqX5I9XxiKAkx3KQpCLHvrTYxIDcg/kVRc1pYoHi+rTw/ItTeDdWefJ2xOtUTk
lni5ZZsVtsDkmEZXiROZfW+2Hjawfo/vGH1Hm3SgsQRO79qM0t+Y8CoEzvQY4d9L
vm83KeYoQdyp9P3+0LiHAfsoob7C6jwndA3X+WpE3QCbPjmR6QLivWsAITH15B9u
7e9IwBoAbUiRBLDzvy4FRREyjIQmq6lyD61h/lqoAVvFDYoToCyp5Q2zvpqLxVAk
Wx6iziNxiZQGmU7K9VpW3WDstyuytjyJnNwTuD9V5pCzOCM9nQVTfCw5OuxStpEL
vaZqF5ld5YMly6fHFEBQ87HOdSJce18miaa4ORVQ/sLhfEZb47oFhRpKgQ1oD1Px
aChw9ab1rYhY6tiUUtfGyWcRW/sUpgn9g3O+51qORZOVpzJwlfcAJrkGllPHdEAy
XZprsqD33gakZ0Uy9Ft0F4qf9xmnclSZv4JIdaij+/A4FFvPtpzJ0kCrkprw2m3a
k4InFH1el7h4c3wJw0m+i1gC3KKEjnbAIrm7PuvEC1gXSKZR656IJdcmCgu9m1d0
DUG2JbptFn2wwvAXQ2dZ70oi3dAfjUtjYAqPBX/D9ZRf50s9R967ojMAlFj6+LkD
PRHNIlP+ys2adK4zpV+4esFqIsvDHi5JZt4QoqAAeOvUs+PmbD4I8a4S8IwWE1gF
k/5VMAYTdTTIH+c6lmsOXnuD/H6uCsYRzFglVtL73+XH6s/8XynHfu4drrF4+Nmj
114KVtddI1PsxkHIatR6SxNwlEFsnOd8eyauStbjMhk3PtzXIf8LA58SveDBV8hY
WzUpWRFH96mPIfVyTPcyuWW4bDaFTHoT0GMgZcFE485zv7QDU2fiU75OomkoAEn+
GvRkxerxFA4Zzlk0pHzK7hLoFnO8/ebFYPl7UV266ZxoZ5pg9J9oJs0noK0+3SxT
QGz0xZdblGQQl+PCAgwONnLK8UuYbyqHtX+Evv+DP1B1Wzebr2JUbLWT7VpM91VZ
HwsZZ1dlFtvUFqqePSbDS2vVtzX2/73jifNXiNoQOyzRYOb+K51FmuMxu1iV7k4b
SfSAxTqITex9iI07rKIsr6868BGM2V6qFkht+K6mZuLbdBKl7bFYu+/13sQC511X
0XYsbfscCwzH2j8xXA4fzj26Don+7ZpuAIC6kHOTAFcD8lu3ltmr83VdaGANk6k0
5FsXR59FszJpmzPnDF5jGDPGsqvkExOQf+Q3UMjmdCB8IJL/P6ZSDeZFKvGD0qn1
36jys+pwFbbCVBrcWlQmj86W+Ua8BJpTBpy93+reahf6Jply+AwZpazv8lLG68ff
0hVQb60o7xqrRHDCM9FxAZJZm2yGtf9SmREJlzrpt/AGxwC76KBuTjuYOP6RKU07
ckX/ydZuoqj7Y8Fo8OY1SSDeMSu2lWrnT5Sd4LnJhoVa3Y61d802bDZucj6xJipD
IeUQx72f4LdeYg1KsfzXzmOu5ELAUlyOlKQkugc194xVPbeRW4Edpkufd7rTOYPe
OGye4lX9yiIylUcnVfdQwK51mBs/QRRxY0JUL5ISOLN+3+QOVpCla4dtgt0BcoWE
mvGoH3pQtHylE0h0NFLqFt80syyjB6qqBOFNhBCIXA5M/F/qM0D275XlRi+EoAVl
iAZVPqrKpNoCuXYAOSVmgdl1G72b6Sw32tE693BBJFT5MJwCZRLQPhEI72uaWitd
4ddZWeBSt1OHdXfSYfrhMjR6wS/oevmoo1xNJvUoHUlan7dE/nFwXRjC/7dB92BP
SsxP5eld11zCsogygT0iwYG48EpAeK1b3ooj7lGADIttOlW9SWmPZ90we8S1TAm4
jk8rdeKeA1QMll8mZDUqVJnZVIR910cDf1+8jdCLi94gkTL573UoAQr4I7JwTOk4
Jg8TEtX8Fy6FhjaYvLzpIzBSeYSbRaifA0+r/XBxzSV3YG157tdunKsJObt+IQ42
3lRBxK2w6vC7ETMII7pmKsY2iCYfLZDDyujdVdjpclQ70wO8l4THqxQymqnUAifj
eK8BDzAdXP/4abSQysHV4awPBzvJDaKl8puFB+CLjhEBqWU5lmObolmcVmyD6wDV
Zp5PKh2SzzNQZa8U5SpDpxItUu1PDEsQjJV14prEveWAcirlj8ftEcKA3yj1wa/s
vHGKNR+4VFWlxAjVIESHb/WkErRYnCYY62BH4JFmxB0zyQJgxmu8AjwEzlzW/r5H
eIcW9/gSjdDEacmDvjIVAGjgV62RX5sR7Ma7dhGqEmsosqyLUl48UDMXl1YxU48l
9Fl1LsaTbxhGSYtkzuI+kKaTOwoEmRdvOwF/lzFKq5BQIn8OINkhOkGhbYFXEYkB
OfNyj48hiN5704SZihIo/0eEzzTXRIcEGgbgbWPrs11u6PETmRLuSMEUIB4GPS51
I0Y0J2Ah1N/akm2b8dNsc7tA3Vu5owlz7VFMJMWDTE6mJMtnRdaPA3JZ0zmiUEQs
vzu+5PiE7VB9i+msaL2rYB4iRX69KLLZePXo03rvF0u2LwJvSp0TvTAcxIUdas2+
qzZ3XxKR8CWpkFJqY35mgKob6emulfJ0zZKNw9SsSkKlmRct5c/lGzLPNaiM+S3s
K+BnOdxTxQZDFTMj0TIFJaDLX4bEv0QHRrTljDk7SMsMoazZGWtImahqpGRiYGkG
AxaTkNukiM/L+hK42Gkz+ZNKgtPHv15wzHfHYokBlLLeSA8hxSX+HrzxKbFlZzBk
7x8ElfySR+Vwm4F87ifY58tE9tv9TQ8m2E3qL7ySBxP0KEF39svaPcVg/brGN8zi
r8b+F3YOgHvQ3bmuN3aSTQsyyFUwsF5BNThgKb7X5jyp1xXj8aAaPnS+A74vYOWB
HnTewqH9SRMQqM0mFrU/0d2BA5lMGt6fqEbgSwXsXIEyu7+yhEkh372pHxZd8LEd
hWXKgUVPGzDgqzMK+sAK0tqQv+laKHo7x2t8k4b4M9LNImJywjr8S+egA86ia2CT
X1xvluC0FId7RTblWVDEmyWM78k+NtisgRg3JeRPRrtUaufcQW2DLhBNUkJrjxgp
IbEkqU+u56dSnOHY2uMI0Mj/N/hDbqkt3D9aLJfk9eFhHItszIIft/XYnjEjJnaR
xeiGacBKG4P8iZZO6T6aUsmWjPHGig246gjvn1TWchcarOK3Nz92050fVRHCg4QG
Ys3rMH5pLywdP/i+sKsaIcfmPRQUZ9390xDlsTP4lbVq+Q1UWzkSAf2qRrCHL2fy
Ukatstz8+v8QN5HCp3UvEa8X1nxiIn+UXVZ+vc1ZE2U5U+/pzA1URDYoAUHo6iyt
GMeN4+AIpDnVkatZS9/7//QPLQrlmuFkHBLyaY1bH99IxSoZJ3JPNGgsve0V7nY2
BwkBGN4nNKRvG0TuuhNDcalqgrVfJY3HEm6ngFVk/n4b6uUVdSxNvkeBuzm4i9Bc
RSp3M9z+FRsg6lCn/kOzFjhF8GtxLaHPmynKuHqIwHRcThMPwNISbStyyKz7/yy+
F8E0dTysj+WmtopgpwhrA86FDCxfqgEZFtTx1kRwJNFcVEnTg962dmylpECJw220
d0lRn5ChQGvuLpLSOAPAesC1hjBhPsgkQctT1H/pJoeIKq0MNo132IkYpkpsqpNd
BJX1sAUTbXRAH0wTNYTpTske01pWWFj58F8USAgTU51AztHmIiP4lTLy+mSo9f9S
dS8V2wrdtXeJ5hMC/0RGOoWgb+fK6LYDQKAKVOjJmx5iGyGMNZXy0rho9oRxcqod
nL3OX5PCSFdaMLyBVAziyUiyFC368RjDFRhRum6z85SplVzEi7CgOW+Tgyx1+MDF
JT8xBRLucn7o5/e0S4a5OJCv18flKIGW06EeWTlCRXXrNasIvvgw6BGpuicBTkHJ
RWYXJKKwBiPu9P/Q6UdquQTFKyaQuRKzLmnJzPy82wqal8OawbXep0NXAFvjKl8H
VTtkzUONT3b8yVX1o3+38qY0cVw1iS1cKU7j+Bo1oVOMa9u59phq2Vg5jS807Wwn
X4mJS/2m9xPX29+0GyoYFfjLT+W7aj6bdrnL6cuSPfzkIENPIUK99/gfAhC21Nu9
3zzdhLSFi76KcKRujE7VRs1xJD7zlMd/cdVUPZhMwIcyD2k0YlTtTu8axSuYPGJO
/9Q7UiRP37QHvfXhUBhElTnY9hR5oT+9pYTe9yPiTIvueOw6tGqVlj2znkFNxrzo
sgWHGMZ1KNSUhtTfMcNZaZCmkrODVI1Y/hcDAEz1ckMrm80ZTIJ3Lhx1c9/2YFJe
Omg82qWN+6frSZVdndjlCSb0OYB+TF7729LT4YjcVdQkJJyq8UuxOPaLVmH/xs+v
7+2StFEguCn/nHzJkVjWEFwU6m6m3T545H8YWE3Zx602DWhYv3CwQGekPu+zFwNV
6/ut9nZb+E+Lf9t6ky2C/aU2+K918V88uTBTLUH6d7py1fSWZymfUpGuy69QaR1b
n8MJtZpu5HjGmKYegNwJ4jmebxYyMFQ9/wUsgvjiN/VSvBhRi8qc9ugiTtW4+pZv
FipKrMYIgmi8yfkw3pKjGvw6aCRnhJvTbSnHvv1cp4Fzps0/qpsw69cAC+9RnOkF
Kzptf317Iyb8YQUoTFyuNt+Ow+O+kjiOX6B1A2YiFdRr1Mh1DY4eC1/3UKRiVFQe
FscZprB6VBLEFH9gala3JhjoZJ5MKOehoaTDfXccTC5zB7/VLHxf4W0ytj8/T63I
tbCPz9qw/7jHpCPGzXIs7L99CRCDaKEnfO7netWyty0GlzoXucpxQBepZhUqW6zb
TtWBGNnAmKqR6kMGb6xPMX/3atioCTAjW5Gm6Q7VvsCujwjsJgIbwuB66pqgSb8A
gbssxLtAd52cgGCv6LftbUD/Fn5zYWHcY9d6CAeglpT97vlNqKI+yX4wuXM7CDWQ
f67Aa7vaKPkBsmtLOAdtAl3mx4xaQodLXxvmyF1w9XTIoiy5TJyv+Kczq2KDmiZL
YfAI7mIKvLCqwTigrhv8As5t68vlatg8oxO+1pN4MyL3fWcFEAq2LmztKCZi3ISF
LU8c8Sn+WspM+aGUpibLRH6BTgtZsD5I9UuAXs3SE/hPHbIImRxFcOOVFeJ7em8K
A/2xzSx/fPlWqr4JpuqqF4IivwHQQjhaKsh/JILkuo9ZZ4oYXmUzQ09rRckguR6x
x3zJOcZ44OajWz0SnT0weWxjzG7813st51Pa2f7qRWUw/p/3yCbxVSOqznpXLT8c
9tcUAkjsGOKp8vFbGczPRmM1DkHk2TyQy/MQz22m96lQmIPiDyaXIICc+Re+V/xD
t0NyKI5V4layV0hVMdGClp2a0lLvFusseHnjPnq3wofbA9vuH0BzN1ZlPzl7VFP3
rf6ZH7kcKWfRdEr1ACxtxXhbeMQPdBqSgfezBFmsyeGkq3HHKIbS9K7E3uoP4/39
gHpc23BCqoYvSFDDAP4I9Sgww6neiAncS1rYY8uV0uVnqAsDmXGzzerfE+tcLvxf
pYyye5jHc1hTJkM3u7CrTRtTvKIlO/5QlZrF+TEbJ2Yc2mbToi2vxKzi/AOJ5aUk
haGvC+G3PWh7AhJ7Hr/3edZQfqWBlOdAID6FWOqkVvOAbPXGulAMUvyz3zj4AQ20
68uq5mFgRYXI0BhgBois1r5OvvnMCCy1BJF2TsH9IPL5F0aI5DsqlJUTIxWWAQNe
IIfK38ND6Fj73nltOzWK7QUGg7BN4hYcnJyq/xtoa347d1kb9HHnfgf7M0SoYmsN
DNWazWzd+GaprcvipEWtfdV3xxawSMaGPWV4TdBoTizM/sX73a/szCezoZM6Eebo
NIeUIQdAF6HQ+Hr+S5xzuCifNKIhDowpgFWKY0IpE0AAQC1sfsHa5IVs/xIET4Jw
+1CWqGs3XuC4SWawn9zfTo/Kgq2W6pMEzWtmWUcsfZKANPe/0xNNzvDbrNemhaLM
00lGADkC8dpxgUj/DQFmWr4ZgKYCtxrz2OT059I+/Hn+fzRmR+3Dse2TO09etOCd
aPAewMt/afFb7rjij1csKWAjxXZ4Inj/Ey2iMdI+Bpncqocfg4/8oKGlARksrC/n
uhje7FvWUY0nEWKW5ZI02PUPD3DEcx9DUq6G35cAT/32DiG8qIGarFKAWXnQuvMw
P3xmARprlKu1AfGoP5BwxKl1wVM4cT/4ZqPrnEVImq4nnTsR56rqSxraqg/nhjxR
Pmkc0Bbw11VDBsks2j/PugPMn5DeLU5nju+clCxyOQMiwlFGvyrzpjZ+kejrJglV
yrjiUaOkIMYCrBsCHoN2qlZzuCYkzoQU2igiMaFeujSS3z40MQPvEF5ZPX/3oxIQ
5R+P02AbArO+QX5OoYzsLioDZZkJv9cqRLF4yHA3tB0br3Q9pqojZ50uouqrgcVb
+38jN5kW5iHEAF0Ak0aJEObWP6EJ3rYiLm74yPOCqY4RPkDhGUDSmWQpeB7cwsEf
dlKO559B4inozMvIn77douxCQDoD0r2JneCtWApUqI1w1f54YInPgmjMA1exEyoC
cYozrOl5nt9OJ40u/6FGnaDhOeHoWYOSj8Kwj2nB4N82EvPMSaH0vHhB1Ay3CJuv
vg+v/dEue4D/rU9fxwFM67rKXT6/Fc31S20SxP5pV+0X9wkAGJ/GC3TvKaVupJTK
RjMpn167dlcGSmgecc4d8+VJRymT1j7PfFkxMxsQUkV5fYF51DGB+8ElGRxOv1FU
Gup14X2RED8E9WsMifoolXnK0yF+ullQqahpN8vfT4uueMQXcwXgH0ixbbiV9tcB
GSf6/WPjhA/T/8givBycMexqoxzfwdIusvHlvWn3pt2lGZoorld1I14ApUQZ4nHm
iWFPTE/0UoKcBG2bjZdvYMbN1AA7j8lXGbHS2SufEWLc9YTbBhcwbxSgTvi5IclJ
DvJHIyeA+43W8ALpiGpwsfS1O7asoXRz72ylaZZkoCh30ZBQAmbIkkjNrYoZWNl+
3BKVgCDGYanwCFWgzjO3Cw1Pq+KeY+5vioVMe8NXrF0vshr/7h7GLXTgvkgvTqF2
jGb60ViJAB7/7XZy5Z7vhdpWeUSFhnhapeIbaciXmLnhKDmStOxcMBh1jr3r/6w2
lb7MNBSC96dQX8j0iyqwtm82Y3lma0L+BpnndwAKze7qR8ZLea8KZaAvtNTnP3OI
Kpdq73gElGcpqb3Rim7F7Olp2HdswCnMuXY2/qVFTXfcZQXaUqF5qnjTW7xWRcs8
9WTf5ggWCFe2aBeMjCt43po9IWaKd4kHjbpUdqvsLSh9myRXyuvbGIrklenvnGnU
mPtgGz5o+Jew7lWsSbcKRbF9M4KKkgjzpxSewe29svH9z129RG88Sc2AsBrdVFm2
b3g1GXOTsgCXA0H0Afzg/CZHf6klydzpn1TAvrkpibdB+b/8igJGtAFFQol9cc9G
VLn6jr/AUGdDVO9PklOmrTxboVXqCdmp8wQH+AkE5yWSzPw5CYNEDk3ojI0e0ZgM
Litmvz61nNCjMqTVaRgEVlpQzH12vzcNHYA9t3qIaaq5GVRZFVjndp7gVl3q0QFk
H/rOrOsLCsuYjCzsH1vs9t91JFWjJfFVR1h1gGii3715mw+4004lDROUu3Pglp+j
CD2sMxqiVf0Ys2WvYmX0o6WdWBQyyTLz3uDCrMu0QGIDNf5GJyMd7RRcgkalEpJt
iT9OIT44bNSAODEmhpk0Dgnmop+/7THoe8/niApQ69Bw7XbbtVSdUCZR+TRqqU4i
JglfYE8AXdQ/G+bO1+ona1owYyyNFLnNyIfKJhUvv/iGhHZjUgeSVlWIKqx6cssv
qhAqfwvjjJd+KuNYm+j95YQBMtfsHRi7vIy2zMJFNJ/dTbNnI7jsFt96Qx+Crq5M
XU1F8tA10gJYEAWS01NtSYGE8di+FLp4BYWChYFa5tUHO3NC1Z0ECDa1gx866ptG
iURPv1QjYcV1kcrrRdk6qaQEAZ/zf7VypZmgpNBVk0cYYQMDTdj7UCKnNWqMaDu8
ShRTn1OeD4eHTstsoGLGpcDYSTb1nyBU0RdcE5u1NAIbg/yAk7BQMymgZ6n8NcRn
jfLYUi6UE/KKh4Ld+Ss3kW60e5EUnMM/VUOjwLycJOzJ1R86AkaQdvYSoFYTsCOX
TQYxaNdwrsD6BExaVDXDVtdVXJKXI4Jqo51U7bkELDAkg1vwSXgUMFzRkcJrFAvt
qtcA6IlyXHR2pUQtEAhOyDSLnDy6XbJPYwobXZgGhzVCDUxvxQzQ9NqoD5V5/p9P
ozmzFsJ2SD8yG0OLIOvEnzaaFWZUetTAIdCM/KgBrkvqxob47iV2MN9PcJLE0nkv
MRxBb/LT8hgWH4HDdbJpIniD16WCHZpiSeZctH2MEn+CGXqKwafkE9/PuzUjrJFF
vsRV6NIJpCMWXxlddOOTgp2TlhkHDQR4cJqTvfLM6QuPvvupwUWxPOB2sxdSjl7a
4RpuMWjlYBAjbX7PMWNvOogl2LI/ilhP3t+F1IZLXl/sBYgqtfbQb9WDD26qxoMB
fScoHPxwrVWYKd/EajRr6HDjF7Dmuyu8dZFh+xakc1ODKeRYGJHUUbM8+xR7fmBK
sXT+xjVexk7HAgFvfdC/T/3Xt99HFMhBS7q+nXLJvn60Gh+gsP+meD219CCpeJGa
/VsjeCeSF8FJJmVwEb19j4tltdItw8T1Ks4r4R8DE96q5kiCjB3AVioGoCHt9fPA
D5mSlyrgV3K8VXw2i1QVjBqO3le/Uni97NAa3cPw99G3Gj7OHJUrj/xFKIBAaxlU
COSC9jW2or6BvPuG8cJdKMlfijVcULDSEmeA1I93+/GaQer/khRe9PdrOi2O+9LB
vF710HVBRQB+4STtTT7/vISeR2II6/ds7gV7BdRpY9FO2DXfgmi4r6VcFXsFpzp9
JHqJ/8cm2+2GJ3rlzxMqAekfeiws4tZ+bVOChvj8YLMeFJYe1qDg93X9Q/zOyWv1
BOFqe+OTa5vOe4ykO5kiH51Zn4o4lIf5FAq5dwxBN5slR16/D8byreTbZXxMJ2xR
3/+a7nQauI5NpRjtVgNarTKVFbojY6rbUI4MKEnPDFwdO3hwP7j+A6zMs/vdg0Sh
kaWdsHaaLmrPwvSKwB71uE0vSXgBwYX06wpc4InSyQZNC0VHnNEeb0BhX2OCGfgj
06tWFxw5Lo0UUVXIKGFVb8nmNFcypi+yJtundc7SvLKuox/FSYrblGSjaPmuyv1Y
M4OQuZSoitJ2KqwakHHkJGJlnS8XC2ZQTU5DtlIu+nGkd5p3LJu/d/1FPco4IVF2
f/jaTKDeGNbPv+P0TyNKylq5+ZJdjJ3chTQOsD3jai3Kp1fbLh9hoxL/HkvjXDzY
ZbuWEtuE7zEgKAIp5xP5nYh7RkLhFD6LToNIm3Hd4k6qFDI1DEC7UJO5Q7cIcKUh
ewaHcEHAZrH88Zxww8V01nQFQ/mxDHG7maSikNrxDuiQefK5XN4OHbrr5lBpgTWk
tVfgXf/Ru49FhGJ5Q8tR2iTtpAvQkBaxghl5hEYkaQ3jyFg/EEkuSvOgiTic1jh7
jeh8oW04BpLNPFu+7YdOAWheSCdaw9wa8hmhKd2j9pFwvxh0xEv42AKAq+d5zsxQ
j2RKWdZJbJZMaBK3nKF9mJ5VaRRx6khV8kCvIm0OqoTbsJBCxUtY15hQJKJlvQpP
O6hvfpXjr1x5JQowyWOvDMFOFm/z/oUXzXfsqz7FNW3tjGN8mBiW32wMTgUukLg+
GlKoGX3lMvtNyWpFpXAbB2dL5ICaqOSf2HRsP42sJLwh7MyY8r+9Dg0Sx5GM8iuk
T2c+uHP8SoT7/e9IxDlras4NJbzeK5NsbScq2JSC/0+ypkfSD3L5hvSKJhSb9dYg
kP/Bg+WDotcsV6qc24IpWLizgtF6YyestRtM4S6cRSeML93gRmyZA1LF4k7XgMF5
WO+wklL/pHByJEkLfXvCI9UgwXTn9UZpYQM9RWrrKSxH5sCs5HC+mfzQlyz/5amX
CGHkf99S/yUbfo6hMoqP2YbY/SFG9MiHV7ozKqicmM4VqT8e1W3eZQu617UhJWu2
n8/CoyCnI8BfMo16BlaH6aU8GY6ahT/rsiyBEriY2kTsng59TBhJbPJEnGS4JtYZ
jGmtbBds9vzqQL00i1JLdxLDXFrl8+5sygWCik6BwY43DHLnupUC83O0CbDkiSwR
xZdtZtIwQH9X6rPxAlKBH0RWhDlu1xEKWtQHqAW8/y3DVhFbiKXX7aQRV5+ZdvBR
aZFsRVXdKjJqu0mZJXdsfJuNNFXvOSe0cd7IrtT+jDW1aNCg7lbPvL732Sw9khcG
GyPJxeT75jrA6Iq7GVRi2scwpsMXuiMXZ04l9x+C0pkcipGAkka/u6mXsSyaTcNo
Bugg3FD0L8oAqaRHZSDsnj+3z2GwwOQw+0EKPGuf3XmrfKznyXwJHa/KwRqQ32gO
QWV2a2O4w+mJw5S4y7Mgvk7nFSYxQnOoc+cizIXEeU9pwgbxVcQRrf71KM4RuCyw
a5h7J3I6dnj5rjYlm8v8eXYR42xmc9ac1qXUvZW5QTQVMGJxTaE5re5Y5cS4iIOr
R10awFnJJPCQR5bTShRweSUJBV3sm2HKYNvVbJEWTPe+iONYBKiSfxieCqkuzz6X
6HMY3r4puS1gKnY12ZA/U0HzCJ4/sW/LTT42KO/okSb0oGxtacaeeI3Ba2UlqL1k
jK5ppYAtkRVY/Yd+3rswjnSHD+1/eXaCEpw2QgQC2xyDy6CxAZNITT2C/m09X/os
SOGEYSzsIOCQG98xLltDuGOtVJ+QeDdlWNOixYO2R5a1ga8RQjF7G2LNY1PwaIxa
WKldL93XxJdE2KctmFAQTpCAQSbdQL2jeLnDShQRrfWVq0HnIJPdn18RtSgSOI0K
IzdUEGZTNng26NQIOKjV0zr3l0skJzvyxObX6v1YwMAYMLeEuqROfv7FtOh3NjBn
2TEKMOthB6jiJdevrfDlypF1d3EzxYV55Hhy5gHYzgep9ziLFz7taHjjSabZgMkk
XZDk4nGAxKd0+UKtqJ3A6lQag8AvUBr1s/CW9PwEWJWk6SNGip7TW13EzN6ufSEg
qhaqdMuKQsx6D9xxY7RXfF2ZI9R1CBpnjJiCaprLit/WZbUn2OBqZFo9PrrzYJGO
fQQl8f5iXS5+7+g1raRMAPsZiCUWJZG5KzFZrGkquO1Eg5TOLgpMUTPsNrPFY4Y0
le0tht6sU1XybzSqre/Xo76tu8Fp/lYN0D8jBdNG6nzg039rxYWM3X5C/xsQZf7T
nImc0cXYVoraWK60YkFdxIj2j9GeQY60T1bi0NhL3sI7lFdgSc5kpt2oKVrMxV+s
dWUcgCkbhzeU46hTTmn8FX4ZBcSKoIrsXmjeZR51Ept1LhkjTy6uoSAIfMoxxOPV
T7MhYAF2B8G5wImus+TIeL1WW0Ezq+0JMesTSWV35gkmK+Wx0UBTcKby1z2QG1B0
YXjd26KUyaCXpjcBGoXfQNYNxCUSqJQxTRja4/Y3KKFvB4Q28mnNAGsJsL5HwQ2T
JipX04teJ6uFMmeysuBz+8l7hcdldFYDwtP48ph4qkg/SpDmIx1+ApvI+OQw53ng
7qasTqionYZVHUlt8JwWayVXm7cS6vZyE9R3CfkIDSArdnN6V8E2yWM4SyXGrYk+
qoaBnINQRiym+PO2qKC+IK2TJ7m4Jz7j7zygWka3cSRLB0tRR+c8cJH/8+6g7S8H
R/aYHqoYkMYwBlcRdqOu31RGTJx6Zs+fawYoyRJ+nKQwt2DkRaSzMvNnk1U4UNqn
g5Qbo66QViVMeiTAq0svfoDP7EBy3vPneYRqZgT3OKFwN4znIVOzoI8zyZXETg/3
xthFasp+NDoJGWv2AHkW/RmLg+0cNiy3JIchMCkS2ACjRm7XJYVjZypZ1Pt3lBzD
CWDfYeN/IrRPBhboTjmX8mcnt+iGTuqZ/pAGSPsL3yrUThwPDMUkeHJRTOkTrf8o
ZKUHjIiw5+428BRWe2CSyVwsoqT2NPjiegDQYcaJFw/e9HLSqkmHsUrIlSbd/dth
CymacWD2VvcUYk/VbmijTtZN4izVzi4Y26QJEG6HEm2EiQSQ2cUiVOUXCtQ5N7uQ
t7MCfJszTLHAqSFq5uF19vQylxRxidtzHkpw/DOEFFHb4M+NB5GthDNyep9jstEO
+5SOlT+qx6sKiWjJgYp2fautTBb+JQUB3qnlvo/fty42hhpTo6hxW6Y5Hns4DK0l
W5dWyyA0wRT1vn9FXyviPBQF2+B5/I0cd/UPyHtQwiCmCwAo4FNaXOarqprODXV6
2rZLFRU7fJPkFJooIUAwMVwbB551FGz9tbgLGB4sZd86uiwoLGTTYFjBF1G5je34
WoXCfwvS2lO9+oGevHYRvej/BuoP45Wiy0qdBJTzOH16IJ349Ve3pvf3MO0QtWRs
VMgkm/F9YweCUHxDVPZlSya4Tx+A27SD374KBP38yBdTYAtr37z6RDZSDi/rqZvQ
cgWNASx8rfxrLWpFO5AAMIhclen+Rv92L82PcYbO++tn8fVFbrZ2yNG9rlp2fYuM
3SiDu6+l+RJU13cHkfhZbkftGVhfoVw3vudttiA68htEZVO6APjJ+NAy7dia+yKq
lrwKdWLnR75gwwDV7Fo9+qhZnXpisiQzRJA2VO5s6VoUkHSHh0aOpPui+gpTORqo
iRBiLa/hgwNVi+L6naUz7k1XeIjU/UYtITytJRBHcdrkN3H8S9JPGOr9NO7D+k8i
VaaTUx15bk332mc81HvaglDcM0AhOvPH3s/7xuJ+HUdaglT1mEMk1Z6A4hJze3mz
Abq/38dEXyYSVsPko7PLtL8AfUhwIBZwqW+LEaqbB8QgLsD84fCx5x6+yHwbarK2
uLxxc2f4CY+qWaCQoQaFU+NatjXGVR5tKnaMCOD1Z7jXbD+MfU3AYA8WCfzhCRDw
Ukxy5l1FUU9ZTDwQXKeDMHYE3h/3Fer97MicnncKVCtbG+gjHAWaTsAqj9Kahl3U
0zp/J/JhehGHV3vSzBV2dV74h+QRH+0a/nTq6ZrXuRyfJjC1h/t1d6BdNk6EjyE0
ts2LTDvnREU+/5TSi4M6+Ll14LaEUlRCcERykZphNjhFme9jV8aeMSi3Fc7rrFIG
9AnCy46ncowgvkemdw+6eb6LyaP2Gb0y83cWT1ABB+n26X7vEIx+Hx4JmVuRIzxE
z6MuaDestzfH1a2yhLTJnq3Kc3Bz20Wa6I6wkY6RRjU10p8znCYaFdAjtuDqmmAj
41jpFwgl4TdIXKmPbi1tRGWo2PxIzrEn0jtYjuK76Ko1oTQ7+cOOV6Jn/CicM/Rb
t1/W/Y2uLIIhXkREm4FmWnYz5NK58Gv5EeAPLn85+epGt/9id5gmLhRbiA+HgaLk
XV5TCCKzfdLnv5h0TQfu5VLJkz4HAneK7HVZhb67zmFp+Xi8M0l4ix9bjt23hyQE
tqpLfz7mJgICAXrBfVKd3xtH6X1TGW0eCfm8ZYizStmeGqAAEafrKyVMen/puJxP
Mpbx/8GRhzeYWxZuhMdQM7j8AL5oMk53B06oJ8KgK1uL64tvE/PPcz562SbtboLg
vwfbpv5CZl56vch5dy08Ujc9mLxYJYTQeflNtJ9hsF7rgI7n+vJqBG2KZZt9gEEG
qO8mNZY3VbBKXt8CN5i/1w2Y7T7eCxom4remWU8FknVLcZf/VmrLmCd1Ozc/x1p+
BR8ZVdxVRacQBXiAtr7r+UuiW1Wj5sepJ/H2lnEkFiaGUfXAqVl3NbmqLlfM2D3p
mQ/oBtanVWR6rxatmZ5tje2Vt/pVI8zxHBSqbVbtJ1X01WEgrFN1mvemDYskBGca
fk4uQX6ehQolVkaVD6BbqvCdVpvS47Et9UN1/aCYJEfDH7RVsXQZFNPNpEW457AW
VlHfRe6VurljaUl3W4mDJcOHTF/w2UZIg0gymmQiqqQLzetuDkPfSMNOxoVDu++D
ZwcW1fBDjSh8yqec6dvowchp4ZNyaQw5v3riuAKjPS1T675Q3rsRivMHPyjRPIXq
t9qt3QiQhS8I2SKpQGpHpw==
`pragma protect end_protected

// Copyright (C) 2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std
// ALTERA_TIMESTAMP:Thu Sep 13 06:32:40 PDT 2018
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
YVfhvaAppEW0qYWodTaO0clGPZA0Cq5gEKHgGgQJjRpcVLCXVSAXZlb70kYjAAGH
CI+ITNgE0i6vftUMLvLzJ/ORnA3QiNv28UwCbB9SBIOYLnVaUBBBeM6VBh8azb+e
QDrpH/QMOvLyAiZdnvukTaSiOLuH35NphTv+OiKZTbM=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 11632)
qfg2dXFNi4krD4wH55r0rmZOVLoufgS9udmish6f/GxF7kL+H+v8E1FztIC066hU
mZFdIhkW1EjY3mD97ZbBIu6yTCgLl/HNpRZLEgEgwmV4plKK0tGsr4b+TDnjJfoq
YYq+3bRcsZRF++4ZYKy8XNzLMYmkVYcT4Ezoy74DZQkFKtMZU1qDYMzoDSlqgrrq
T0r2+8J2prylQa8XBQENVygbfKONpfem8hj8/p4pKmtjlwUHQS7o9ld2xoomouWo
s08leZadIbV2w0A+OT6jZnip7sqDorZewmjzk7sNtG+YUYyYoRbH4YahGsDShBkn
PGZdVKAwb9oSQ5wA1vI5aVBu8uHcqvtomeRMPkHJtk2UvDNIHDys+JydzmOOuUD8
lYIPlh0rLoIYbUltI5H4Qb/ELP5hdiCfAbQLcPtqqcnetaOZ0+HiC/Is/qEHMaHM
ZoWF0xbILV5Fo8wwbg5Z/GXmVVeYDsLWAyjk3k6wZUIV63Nw9cKXzUYyueWZcTdB
AN2r7/a7W7ung3V9RqAOTh4jKrtnXrdwJQgR7IOBaabuTfGuZY7DW0xT9wSNKMcO
50MDPNlmwYBoXgyNM8Xt+mTCXtqDYRLi3SWcXI6A12m423HGu8uc2J/+TtlRMOsX
aPKNOieHDWuhdqEk8BmXPA+tbHMc6E5wDvIKvxAEuQW+4ey1C/rPZy3a1GFtkikP
6WlPFzCBZ4f6mALUpTVZA84rdY/doxt7KJ5dxZZER/p0WMusHUMCIJT3SsdXwVcg
mc2hgLLo5dygM72vjr7FPGEhlFbL852zS4qn4Gc538bPcKBT4U+Qxj4UmY4HuSYL
Dm9RzjBMX7E6PF768Wjx/s57P4sZ4N8UJ0aulVcQXoN5/30YTWzyBtvpgv4ogDmM
i48+3TLsdmdSlFA2YgYjpHXZPBhfMKQbyuYVYJOJTwcVZkYlF/jcZ7a1XsXICJez
E6GI+N0pEgssOZtCFIERFUVQItmLibjDmpBKM1FBpMcu0WY6mIo9OG335eTJDJn+
SqV5PlizA4r4QSVAyPjPvhUDfkLZVI+K/uFj1w/VQm/Nn2/jbjU0W6k9OUpZRQkZ
T0Cgq2S1N+qdnGEpyEHNsxR1DcvmnZ82VoVGLDIHejLAtYmQ/aeFeEGkqoSgZR0T
CwBZp8ViSzes6tzmeI/CDXwReO+CWNOVZk10P7gM5TRqTiPaFdPnJxzALV7jayqF
uUE8dPWdCmtV2Mi6ZMa3FUJW7Cn5BaMfHlm3JbLJGsYpqfbtheuQdpK3K8nBi65z
9TCjAquGdR+KmuwqWeaL20PCbCG7PwflLTFCJA6fzPCd0HHwSspKQE8HxT5y1Phz
6sRNGT8LoJzvoPIv+MPFKaKAcMVcYm57rAO8qCDmjIaWqe4c/zoPTD9bYdAnh4Kk
NI5P3vAWOxLOW/gJ1DuQpZe9LQvuPi7GpPMGyiW2VPnDACrNXgWnLSZOSHBCM5P8
aoXPd7Yk09vUA2YJQsUJ5eJqEv13QZmOo7arcBs4AsgTcwZdaIPEl9jvff1aIB5N
1pJX13HB3zersqYL5xLtaOi/Xg2jWLv/Nm0vViVDmHkIkHfJuFRbu5Dxhly92xKB
0Vh2c6rFMsXNMSH1iQDxCDZA3jmGrbUyWqpjAE+Rx92JcZJP9/+/33jFlqfSzEqD
Y4cbEblf7BCcup6MuBVWmJW4fTlvlbQD/AiHs/YmulnPdrzN9sUj6mAEzXALrlgV
9gUtsM8VYwI0VrzwdSn3Cl117utoextSPJBlBiAx46KycbxpucwRhYYjcuUwUBY0
horLPEIBmnnx7vQ6hJwcNndurbqCIRCY6n+lLv7b0lj6LFu/N+A0ztBE0Ta+nnfd
dlo0CE3Z6ywX7+uBWJa1YeNYBq7LRF0ndmVdXEaiwcIRVs5f4QB1RDUvgviVjQsf
QWVOi/LDiPXzACcqwBicM2omjKkOM4KCT3Y6g1rT4g5KbGDFUSLITO1QSWJCCp2p
tSY/aakot21niiVFuGXCCWM1pa9icj+n90wyms0ZPIdGhuq02INg7gfPeYlTL3h9
9tz6zxlT228RXNJEQ5Y7yk2Zc78hXSPiPq3ut8EzpFGaFbFnle9hUGKDScdX9HTh
9Bw3i1v5avDN/Azo7M/ruygOcg4pucdNH2NfI5iNsB4fccfAH3+y0xjb7Aj//iQy
FAc0FvR++HBQB3SJeoJcf/v9XaGPevLOi9XfYiYnectWr/KUHjGwXbgJtMlxBDPn
D5s7YeNVaHterYxF0p0CEOGriQdeud3N5VUma6l4ov52u6ozcHbeads3GJXK/hfj
7E6suQb0VqYo3j2AW63LhebRNNM9J/Y5tOMRq6gqXm7MI4Fo7nK5ODyZKmd21/IF
/e/SifF2Edc+IJqmcFeLx4PTgPKjpsZKsd5L7c6ah1hKV1iijPdsoekAxwD3Vy0e
LHSvvqvZigDOAZqv1yUZ6tjZK9wTtVGZmx0+DkK33wPU/682f4TH6ulj4u/4DIMr
rxZAnXyLv7mWcLTGrn6PZTQoU/pFsGTi1KSPpZs5SUmz94EanonO9BORf49u2Npk
1+7rY7O5d428qlO40Ntwibm1ANUYFmfACoYN5DU6hFUTs4JaVjFQB+G10wdrOPYT
s6GPWaVP3KqaIqqhYiNIhVCPJfEVQqc84sGnVHqznET/wGOJyEkGhuBYdgvZLLHk
3gPdsAO4YP9qcpL5G7GV/ZJTA4jRfB0UrNh6d4xExuCGNXzvbzMSmLfGqHchVp2A
nhbALa8IV+x+FaRBAafAIzCZUIbHQ4nSfOb7N1HQJvIcLVZWIewsCxzwU2T2SMPo
XQhpxHV8uSN1JCDCK8VSWTfCFZybwEEr1Yxp+S22MMRMqhIoxfcCKob7Wt/jh789
xqO61BUhTIlDtBaiWN5aPcaEjT7cZuV1sOV+QRT5XH9EwXg9W9tNZeP5Zv2S1tDI
fJjAoSoINecQlKR88isyiJ9Oy95QCbCwYAsttBy6MDt13sTE2VfG4q9RSi+3Rpoq
1WChNdEFnzHc0VJhlMk3rQIRi1T+BbPLJqQSuHgRCI2NI+czFnmkLlFk3QAr4K1B
vYNbf4SUMM8Px468kLMEFW/MMtXE7QqO+YohFJ4ieWZwEOFviqPy5TQaySOYF6tm
UVUwcO3RAIVJ2ONzDHwz0IvO93EpAvfk8uSmm2cL6pid7/n9r2fFhbpukLNU4b9Q
Qwe0DvYhJ2HAmfyypmR/HQ6zoJD/LtcwvoIw6MNnfrcNelYs3Bm3dsIZxbaDIq/h
jIMioFXU0I9X876S+u4EFP0gkvPyrVQf7CuzAXbhrMvTpI/TNmukOclKDIZ7G0Ck
9l/ieCfZLTx7saN01vgrpt2bUY7ddFJvob/wbDcX19FHLTwir1gvhIQkwh3dChIw
tRAloiNN36DyRkJFmdEHfqlg2Ns/O89tyntsRAvxVZZJxOhorReb4QmdS+gRmwrc
N2EXX5IcdSqftaIVfTnFXPuI9+AzmUW4F21n1Uozy7nGTihRdujoiUBNNLp75iO0
wZWe+L5hC/z7JgqNcAtBMGTnHamddNf+hDdTSES6YC5XluVfUKIw7pfUVyqSa/Y9
f8THOJJfA8Su2xtr0wi+zsldLvbwQ9YIO0pA8A0GHXna76XQ9Zw83grOHrbb9rkR
LWYVhOX36TSx7qyLE6Q3KewQC9AVzEjUka4+WOmJwsbJM5NHiCWKVFEtEPKE1yfM
aTu8LF9OfINlzeUAcoa7dMcYZkj90rFca9ItjTK4DxcRQmC0Rxl3q/0TmMkO9zcD
Wb/cNSp/buDtRTZJUAAoQyoMIQhVxjr05QUm9MryxHm48g2sju5TpML4qdjFUy2x
XGeDDPWLaRmx9nniIqGyLRRUA8+PLgDA+CnnCSJYCPGXYnWDm50ndr++kTPrCDS2
th1WAGeI6GFHF70ad8yAMLvaRHeL04eQbOLocytV0QRFP7RTc8Nem6p0Td2hhA1f
hSLWFp5jlm1hmPZFPG3TrigJtXr2E7OW3iyM+i7o4Se4L0dfq5nwYXRLOhbqFZv4
g/E1tpj6jE/VSVO7HEFeiwsuZpoMljRfpfWdTR/qRsQ4QM+m+3dtE526p/scQzdz
7xYsjxYCP1BQDLlZMydYA57TUetIowI8DIMonDIcwhBew0HymzU5+DhDvGHKUt/4
lRSbBBawVZYMT3mrbUSQLO9UrPRjIYfzlVhgBFF2T3rvnUhNwI0PMvsKHQh9CaS1
EoseJVmmz8SpJMSaRQuZWn/nZfjybSUJjtueh8czPVDCSGS8WFYd511M6vMOmFLz
dE1vlKnVXrMCiwWV3U3mNCUUVhS2mMmAdo6Mtae3F64VVCd2rvyGCNeOEf1zJ3Al
y/kwh6P3M9oiiJ+9W7mHSDgxZ5Dww5mdBStSq1cL9LH9m5Ejacn+Pwq5Ghxp5ucW
4HmqUEgubVnogSfOxln1FpEo+DjpA/5cZL9rfSipcn4SwKUHa+kDk03bifhyySyE
WrNxVpcxquneX/mADQRmyqRXbqvTPdaK6IVAHS+KFT+s61PF88sizrrFdHKzTFR5
gbpLYPlQg6nMghjttjHSQavrahe5dqZgE4ZHanKo+JUVEyuf2djQYnQP+4vVEYMW
8fsTwv3j99nspBLNgYL5metCYjJoYU2GE5uzwmz26wEiAU39aqiShoPh8zT/wqia
sMm2JhZbPQKdZ111YOeORKV+LpwRkBNh7l20WylykqmnNHZNZTG9WLH1iWbGAbxW
ZT8N406tDqstY8gPBVs4KzvDImuz7LKbRXI7kVXE24uyE0of2YLy5SZUTtbi4WCF
zXZdFaiJgQK5BL7UiNHlnyhkwanRtEk/A7R0bHCVJ4BM1MtNTopukWfQEnNtldYW
jhX3R9Zr87BsVfqQwM+WTiftbcdGzqa7k340KcyU5wvPKWzzBxkhRgtdN2EB1HIg
g2Ke1TvBU2W3SVqPAVdMsl88iUaH1IlU/6vg1SUhq0kfKKu95eNIhQsNqNMEBDu2
Kg5ZhP0I1nBbYy9eFfkozcc+733rpFNLE4yyCK8mBT8PVGBXTLdQb8F42H6MpAkk
N7j4KDJEhRSkQYUbbm7L5rfaW9ZsUmCMlt8G5p7PjjVObAMyocZhHMY1m1aKnexi
V4Tz/5yviFkREqdiT/aLIlm7Yculle554lQDW1vYwnKQ/HyaAF4rRNSReJtbDp+O
4TnhtX8+cf9bGlRCGJiD3bkTCMfGbsrVCChg13zxvKHJaO0xB0olBDyL05Ozrv+0
VaSjst1yfU+L6d2ymyNRIxjbAZejuDJoBPs+PmsmrZpvvkNm9cqxDtfrza2HN73l
v2yrgYf53Hald+bGq/Sx3eGqe+c2PEds1K9FhjJHqD0YreQfLn41NZBVqrTk4h63
W5610AFLQmY/ZRYgHs5WWJSfBaGZUWZiISrRcX/sPLJ19XCuvrQX/14KOhKBve/N
q1upCyGq04p71gitS29NEVds04dOFKVyiuAiyvQWFzMjpEvir4bpsJ1uQ6v2ye4B
u7vjSldjxIo9Gd3tHef1CUjqtEzZD4VX7ZfhBFuIG3bKhmNNIT56Wrp7B9Qm0T+H
IfPTi6IfozEQ0UAL4kY/mFLzp9ksvRlj8RFaR/U6WmOydIajaoRBXSa//8bdNqLQ
oc9xodN1y8igEIGi8iCDGP1MNk51HlgfVLhEh9IWMODqnEexXFLHzsbHADVGnizW
lneVvYmyhSgRwsdTxkWTLSRScUdqtMN03fztuH4ZoxB7/uh9jsSt5fUzP1PEDuj5
nQO1Ob6pPeM7NQqVNjEOpz8Cj4cDaqbunlfyeahWebpdXJvqVImqA+F/QnoUJlB4
Y9LVqxrENeuVzPDI0Jh4/EjOL/LdzuZIcQAGvr0lp1FQeSzP/St51Bvj6+EhyTri
hEuG/XdtEnoXLbe9vWkkfBhZEm5UkQ6fq8LcGya3pjnQAUspG4/4D82T8qFh1ToZ
h+LM1CDoJYB0NP7feAjxiPPW8sBeOL6YoydQUXxwQvOTBDiYjqMhOqcUZAMWFxZP
AiTseSGknVanwfVt5NVJApBtIXmR7os1mclTWMmma3H3DgKAeUocDXuV54hueZYH
lRJ3re//CNhJszhoBCLUIrN49mR26C/G/Noev88C7r0GZZNf11+134h0oQxAQJLY
umiSOKA9iDIXbLdrSErWFkW5NOOsz7aTVKpOh+EeSGneZC+VlEWW/y531H/Fc5s1
8SEiDZIzehcNhNy2+P7CoOPWUlHUMd11YmtWDX/9B5UI2mh4ULEEy/k+yfwGau5v
MGbEryokhLVXGhl+54r0hzTOVC3PPT7vTp+GvE9RE5wMkpDcGO/9QjfI6+FCRoAq
2Ne00OdvkNdoQYdacp+Iyoyg5RsSM7uGrbqwW0mhfSDIaUzXiBO+4kOFUycz6nwT
KmtjCYY/9nJ09WXoh1hLXXNCDZYUlc/VHQOf8RWtdSVhYAb8p8AfNjF8vn/BhZqd
L6tTMwotySgyjuHjOemsFrOu41G44z4jdbV+f+IWi2vdHDSxPft1KO2BBo5v81sI
2m0QV9sme5tfWT76SM/gLSjzlocYTkawudGu1RSlBdt/QgcJFuM8ryErI7R8l5jR
IWzjhXHlmjjsNymO5ZidBJ15SwOjR5OqgYgeqxuTV5VlDwlHKWYLTE2viaFfze7s
xGN2cWlxo4ly0BbhTLDLhlG8nmQCZSKLWwFmfs+YDNQqGBBSIJxkgMgAUKyI+3uI
ECYz77CZTjq+m0ohSBbtzaD6wlF1rxe1/qQO2KeCvkmUhZPaC1y6oLxtsjI+LqS1
PehM5NZBf4TQT7NvhtCsWFNpSBm5mW3B/w9rSRW6ZXL88+hvI6dnZ3ZmqCGoEZYb
Xkh1uPCLSb5X9vJ9cLJDMx2kljubOyKJX97Jpmmy/dyn2+Clq0mL2ouUMJoOhAYd
iZThSVbLVJJ8Ffl/ExfXJJXV7JnpbzwdTMWH4zvAtN1fbFZLmcFJxz0JZao+CGv5
lMjjm6/gCTWad3KKSZE5IhNJb4Z51K5d1ws1zNJkjlzqIR1m2tqQZN1NtmeS0sfI
412KLmRqDbmWRVDVhidBZfQuCFQeFgKha9ixUEGPyMQvynsypZawtzOC8fyGyNCe
27E1ZunZPJ3UhGLEjPAJhV4OY+oodhyVvC41XRGMi5Hg1WWs3UADX5pmeNvOmf0i
g7BcoCShCYk0uOPzs6QSkU1gj8lhRkApy2IOiZGStmUpDfm/DU3QWU5AXdz835GJ
2X49vw59Fb9Ibg1XjVxhcSr4XOnVP8bzzVO6mL1jBfiEdLko6k7GC+PS9GR0nw4T
X/0kYYt4Ou0kPyV+W9NOMt8KCUO2oDUd4bTUd5LNXcJHfF/8tM1mTzrQkogYW3zO
NpyDRA2ISXCJD3FSWshUvDPiDjtbaG6XNGu0np81NW3bCzGX1KLUmCSAfjpASZt0
VlIeaXzunOVuhAK/vlUISHz5t3EyoO5p0Vn3ayNANHrdpdOcLGXPVVpsnfHOV0Vy
PUxmq+tslqQJGltwBGEnvFLuF1LLkHGAWbgEvEELg8PHtHgmdNYkvegZkXknhOC6
I3uHZuNwdcbmCFwNdqDdMYQnsbQGeaA3iwdhXgNm4++MfC4gHQDFNVMir3MZo7KH
UjP4RMn3c/ta6zQrbmzUbLCeNFiLtqsiTsQ1K688t/PT5e58CeHelml3Dn5VvI5N
zsUB05WKJDn1K+CMSJ1TriYJQsZ5Nar0giySyWsyIx8MQvHzeyILhD5xZgaNSYxR
Ljnv++VoeDeJ5x4bzpFp9IHcYh822wyQp2ntBpCm/ZVSAU2ZcFwQSkAxAl1Dx6s8
kPzCUifMv3OHwLTHzusHrV/eUudxXqdyMRtEx2LK4t4xDEa0sSeiiVt/XfT4QHmM
rkWP0D0iwYAgb1j6Ryv4KqrNuk+MCdKcEiq+FOdGK97pX7b0JcBOtQmUvTY2cjd5
dRd2H4XB7UjDc+yX17lQ7nVMX4Vss7en7p9CNNYPmp+FjZ6JZG9foCYstWSaBoxU
jeWl4+AKdPAHvEuebqznb1zuO362/M0Z9v09qXr+O1lAXnt0IFPSL2sULyGVplCt
kmAXWq0G3uz2srmKRX8faTToekHfCEOpzf8Upi3MDf+QOQtRZ27NySwJ7z1fzLeU
j3SWVaEKTZHx0QbCMQnP7RHhQsgEWesJbGGmthWtJqyWWV7rPeRNmVtdFcmhFVCG
i6/YaIx/d2RpmYCiumJBVAboqXfmNERkI/RGJxGTevZGM6mbGtA/Ud8lnlNJGX+P
EXBrBhnJyKN4y0LW+Bds+/nlGgjmDI4FTJL9OhFdZSG1o9SHTweHzwrH/G/lOJFT
GWhelkDEevHr0BkQSeDTlwxM5n5wUj/htQRNscmj8BrurKy1IawAQ4p49QxB8EPU
MEOplyi3Wf0uaQyypNb71IRIGdzb+K/vNEInAERJDlJ0EPb5lkTxBZQXDCuvOXM4
YbXK381bHhH2cPFefHu4kAckiW2dinb1KIJtSwc3IM6ixTlEo57+CZlxpAB49DGG
AQMBMhNDkDb9oAD0uS0WnKJ6QDglZyiSWUejzX7Nfipf6Wxht6PjuJW4YnSbn1d6
5KlLOHK8od2YOu+YNW2qzPIrjO8WDnQcexULsPPD2opH1JQL84D9S9fBzGDILapj
wkiCq1SrN4BX+WImkvlzB9Vlsm3Af8kAr242f6bZZSNQeuvV7D85F3iaCPeI6T+1
lix1Qji8u9lwD8+8XGInjozmdp2IgnUQimHrIkoCdFxK8S5X0GD05JyxEliQg1mv
DZVFSMoYMbk4OHDIA2jptdfq+a5V/bA1PhNOTxyLoaDEi3X1Zx2WiLxXmkvi6wd4
CvVwq49OUfwCim3xeDslcVedy46M1zOFGg4C7PBObLvGaWV3vbU7ierlYBzj1rgj
a0PTd84FmEL60SjCHUIFHUQH3zkuqQh6+zT7pAWR3q7U1p8rhq3GvGGPF0Z7nCbM
c/FlhfeY5ZmAN/Z0zCxRLdMpMxkWHuO1t51vVtJCjWFN4TJRYmlKr21ZqTIcde5M
sW5kxcmCkzX3P7Uqw9NjLqRiXtgQnMtPPwgk/5PHswYRQJ+SkF1F6OEofz48OMTJ
O/7dx/xUo5WgM5c7GP6zqq9kaPAccUqkPhLpI0lsA+Ek1N12yhWDiyRSH4YoqEwL
er5nnUgWaImE0gUBvCygyVNqystofAqRohXwFvUGr04zwg/fWtXHLjarbpJJEh03
UGc8ZCOL9VlQ/z9prAbZUwieA19+Wi9NEAMYxTw5dLMwxySaUKvUBpIcJJfl3HoX
7Bs7Zsxf/lwkF/gmietNv8fhuJs/qXdVUvD2Kg5+WbMEgBnEgkApohQmnEYLBckA
EOZUZtEPbNuMKVGlx9wW52/Z5rQ0UROvnqfoVQJP36sa5uMbLrOmKj4EIfApblLp
7QSNPmxAyrHJe5BY7suYQRNQ6UKuzN2hh+dSIEGdNXQ7vMyutJH9Rq8cffXuEEl7
z4KCZ1naWIJZvr7Cde5BB2XfSFmzIhFcffElAbwkYzyWCePu/9jCOd94hmcEMGec
2uefx4ZSS/luZOIUPx2WSTdOad7QEIF576q0b0rJ6fy1x5GmhJzpjo4xl/i7lyC4
PElS99/HPEkK0iaYD9zkOHObcb3RMQFgHG+o+nBgkDAkpaarqDvKoh0uPJ31EK3i
B+QthoJ+11DBToXCv/0vJYxXQMLdK4oweHG7dgUwGOR6v5ah5HTob15rl08elzF1
A6cVekqgsO2s3Yd3u5PaFY3NOr7zQxGawIwgc8bPB22q+mWsjzdDah4KbkUQRJIn
Q0Kxks+bel2PuTDz6QlajRJshh3e18vOxWhl/UAwyNJCEpzoMwPSLeXP7Kv4VLth
mquDwQNzJuxRAXmKauys8QLpYuZeo/0zcscBv7SkQR+iqmEf+Z50IhxVZvoxQ+QK
m0EHuMtAUQLr/n0d/RNvB54p4//PtG9gsTXv2MQwUJksvUV8rXG2yJvXW6bUGF+h
/g0ypS2FEVKgYXlletZAFgviSoJHGSFzxxPfT7ehnpSB5ErM+0S+wUQ/rfD9R9k/
78mdiQi7B3qLaINvW+0aOrb/BR3PAzpQ8wxS6c04aiWQkPf1r2/HCttBj0SiIFjQ
UwGyeLja4077qUT9lFRypLyqSunUwb0ZXpZohiCmKjoCWqurzbDrV2k35z3XZSH6
yJQHVe1GAD0Ie/eMArl3nhmve+mRBLZndGLkjc5/X6xx9NizYf4z+Ua9tjKI7yJQ
d5WhWv7Tuhg5HMXlvpJI4egDnyiHSkc7WkQm5BtlX+xeYWDJMgZ4pksCWWDzH9pc
l16RX4JNBK1dtHXnjGI1RGB/NOGdwqdZMsAUF8H/Lm9hIeXGYslIfXOYoMjE0jss
zeps+XyjulSqQ1Kpgato+OXbRQ+HlxXDBoeP0+3UxwsANSVolbfAPm3k1dAAcz/H
NwtEbHqpzfGoxVpEc56jqLgxOwbfOfrdwa0sw5dS0MmH3q9y0mKzl/FDAv3FmzOo
ijrTZh1m1ea+VLqsNlnzJXYc6Jwc/3ZKsBOqljmV/QFiakwK91xkNY3I42lLHNYi
cFnjNjLEu0d63sPXm3YI2sqSkyzv5XhTiM9FL01+i5xTPBpSzQfZlFP6DrMAklSb
fx4hrjCKWC4mKuVQsiWVNh2zSRXZ8RE4RzTOwp8WTyVSFWhbSOG7DYB7Wa9YQHNL
Gd+b3MHGQHTTDVADhmk4K2hK3IuX3S+KjhcrVJsboi3kIPRaMpjm88ZkiVTWXNvf
x22xBAZzKoJlzls9Agrvyrq4LT600M7pujmgHDHA4xvFgza7zbUbUu45s3Cg+EiJ
ighQx3C3bnL/kVPwuei4Pk0RO8G6zS3hbmVKhDqIvfjpa8opLPVFRdKqrDuusjHr
YusjTsw/thZQMmONQeAO0C65s5ji8krq7u+yBE51Vq76Ne4G8T0ch2xsdhOXBTUG
Q3wtMxI5oPf9jlsebyEO1sbSaKzLcRm6tg3b3h2K49iVU3+pZY+dDk6jGVEbTPI9
mVne23pL/EvbK/edIoaqsp10JhNRtl+snrnk1lr/o9cbEOFphVmRQsOjg4a9RnIX
JvzPcSuvC1kTJIYT7FT2bcYKolelJcqop/dn/bY2qxGNpbmnq0t/DVvt5OugHHWU
Y5IOtucmk0pVL4TsQA8QauceXDA4VfgVTLgABP/g1D1GnJSTcPtcFI1rCrwpGTSG
/oX/qYPoM+gTwYgD10wzBI4zgPheptRjArm1VvMcFvuJecho63OzK5jCFPaY7KhB
w9Jyyh3SviYnqTcn46xkev7KwptbkglcpaTZ5LFmJjpEF2ZtNEORlsPdC6L8C0gn
O63Hz7FkuS/8vw6AEiWbCIvdCWPB+RmcGRdmhOqdvhoyoe67MwEOTkRg4SrWyJBx
gdmtNllZS70SzPCUAjqGjhV6h7Li/iofJmFdSFHXpGhFt2pWA4KBZJsx7ur7tQw9
x5xnzaClJlnYcnmqPbLPZ74PW0AwXLxn9VqJUDDTypse1RjaXveZs7FpTMzq/aUy
04ijZkLm1Z7uyV4WtMYqeQuINJW3ijLMywIg3aeezF4SE0MhcNkBPstqWX/PnW0G
psnzbt9jjMTK/EDV9nEgnK0LFgNM31SiF7xriC9d+5bwUWUFf8xw/LKOTnRVbNux
Nwgko8Vq60rZCprFDn84zd3u19UWGwbBBsZBB7F1Aevf7M7ZNsYhuzwSoCoZ0T3t
Rhh+hShCmqxv2fGOzjtnhiVD4qM3OJYsJm3Ryy74EhVjdi39SpWESLxkH0IwAqGQ
+BBSnsaO5QCsDDDJ1TIViC+6QLjeeDeiC4CJshbUCZWWpxPDfnEIsnCz44LHsDwe
jS4eeaR3JFJHHw0vP9x4bxRZPKu8K0xJKgnR03EKAFlQ0BavM9dWwg4USy46aDqD
cIZtXnKbu4QSTD9b5gRepZOpRc3xSQuFYw79SLXL/vvAU7XwjKgk8Gdc/9DUWD+a
pzm1NVk4wblzc+FEYGVhElodHLg3nS25IKrelqkJkBosimJbrcjnuPP0hCc4qI66
6ECkByV6/QLNiczAwSsW/S8xTlTTOHc3PsznBSj8mdgtmu9vDZRTZIeLvsKBGcce
xQfFw8DGLw8plmKOHZ6xgAjl7s+S5fvPU6zjOEwAnEwCjlIZOMb1DTxmVHGW9BQw
kQXk4tKiOaeud9YZrvL22D3B+vyz32r+Fkxgsds1ktj/SVwqincWpcunNtbhVEQA
CwT7NdPvWxp91WL3/k23qgA6V0aBXkylr2ZsLkq5rrGz6L5ovBnP/zeSs/EZfnn1
qICMOF/07DTSz2QW7sWHtF/RNeFynKMBQvf+0GM7D9D4/wNjw/nfIAfMIrxZLske
Zp+NQm3KvyVvXzfHQUZKPAPg9Gp2vzu/cka/ffJDCzM+9rsnY1+b6fi7hN/OcChH
KTHAI27DvkkQRNuqYj4mo+CzQPak6sVlHrFXT/AJkGdtj4Rb8gmlLuljRGFLT+CC
MnVpyx3skkk+rjzqXUW5PYy7gCmGnC71us+a6n2AXS9OgaPpo3OwuwnoXNiVmN/G
PoI3ueZ5ST9690pQKVvQCioH1AEhCdY/IP2witJ4wnPqyZSvelb55TOINiZTZk1M
mBP6239eYeobmvZQ9D8UyTW/mP/Lyz9WxelkhldrNc2JVsMZhLa46kONiaq3o+x8
pQzF8r+xM1Y6/1qzT45PU4mSIzu9dYCScQhhRLKegkoKMlibTghec1XyqqQltjxe
5WbsoEYfL7PEBuDvCI0cnndXzbo5Hhk8Q3eCHVuvnDuro8CoItk7yi5mjwFvT9V2
6BePL6w4KRXuwwJxiI7XSoWsaEk2abfEA7PeRX0KmJkUx9gqs4K6cQUz5AgOLpDm
HNcoydwOGSFo5OiZwDeVXEXHYm1IPjoQ+lDOHJwJs3FXBOagCaLwqtlqo2XEA/MF
K/QtTmjlzOfCggu8ap8i+dqg3dcfa2jdXD/jdwDvkT/s31DJ1NNS2cGqbX55Fse/
H5RsYrLslk7/0Ccdm6Y6pirjW6YH9wCXHc9lrVWCMuAaI2cefm61IdfXhXQiWM6n
1pdI+Atq0K37hHR2q4geUYrDcYLnH878m4/V9/rBairTHWXWEj16X4pz9OuK9cpM
WZeaPNLHsQiX6JVVYKBpFKpKc3dV9nzdp8cWG6byMlT4Xs5eHJrTNyIwknRCCH6I
5nHI/P/XL37jWko8jP3CW+9LPIoV2xQuR6/zjFrJR8ShWmRiEUngyv/KHzajFsDC
0s7Kh2eLJ1GoLMxVwa7iNPRixhX7qzVG0imvSyFAbBBtRpkf2MpQFkTBKhkh4/Ef
ygn8PpcDoZRKzwlTLE4u3VzX0ek+vvyRgsgN9o5x+upKWpXre2/c8E/CnxgcUcYI
65v2M4FTpsFAeCRWGmDtnWBHEri+AvX9FnCh1cU0IK8JWlwSqS71kk2HaNiSxxRn
Vbsi6Z4MZTSD6xVgr8aOINDpnc/XfwWo8g8b5pQX2d6u/nDgG23WXLREBvVFLkvp
oUW8YV6ndHKN4P2C8B7T2XdqnXN3xw9EB3i9wWdbOZS0Ln1Ipp12pB7KHOTUoRMo
F891lQFWKGnNmNm2HJREcb8m4dZuk01Y2m8XCC9RDeW805qFkMyIf/HHAOyTClNd
1+KP4Ar+ai+mywrtiYYxWLBFDWadWSknC6ta4w9SGYMUk3zQlWGdBX1JBWE4hf4l
/fznfn03zSmb995zXiv7Qip3vlvSSzRkPEo+4w+PBOsQgjBQJl223CdrlSAxbMnw
Av4Hl3K2aQd3nYYZlT3KI7hS1Eo0imfJGkgBfY1IDviCzv0tFj145IWF8ouM+sTO
/I4FkS57ssvYA6bdwW2fD2yO57Wpg4PPOX1B3lKeD8IrtBNEApbAWSoDsSep7fzC
6HSsNLJiBh6NGvISFwEewmp4Fk61GaHjkUTrnOFeBfDvQRpWl72w7CNzPYgS/Oz0
FM6WmVejBtkpdRICRRjwtxHLa63+p7Arjxop9hQ243NziUtswUszw+wJNrImzMBy
vuDoEved58Fnwr429K8vMMmsgJTaIGeJ3OnIFBoxjSpifK3mf9A9yDzGbfUlhVUu
xzxsIKPPQ3C7DPxRmxCahh4gRuqaKtSONSiGuQAmmL8lfKQhXp8T2lWCj59mmWoM
34c0Hyb68rWm+4WWzkLB/53gEWZRm5O/vyqdM0OC8tmX1aK+c/VWp0MX7paXO/2G
Ao+L6vAWeXPWBIeRRca0Dd01zLN8sUYKX4gDqutjpaLz+2+6hylvYh6ftO7gRoAv
tf6GkBuK3C5j8ZJGjexfoVxOg13knXdFyjsrz3EKaIgTORqXeDaPf6GtJ8LmbXf/
+st2D4hBwrAEtt3B97xP5pQW5H0BGXbd306/hMnQleio+1MA81rwyvGww2rBB+hC
RfGMWYLWnAJXsORNnlFoMqdb4TSCV85TDn5vBs03slNZ9fR1D1BAZsiHBx5vB1qS
/dbKLtI+3VyKMHIDTGd3CfEzweFz8BYj8mNvgmL1f8FcZIVjDzvGMTpY0y9MvOgX
g7C+yk6SBR4L5k0zOGUSA4O2qdcNOUpW9+vXdAYpeh7kzPCaGelw2MUUpmNnsDKr
RAT20a/gsY+MJCc13f9bf83bmGCkmAiR7rqVEmcV0X+6AMuu7NbyT9XRZhdqsNZr
H2c1tisPi0uGz6HpOB5FlPW7qo4sVziaRsJHbWhsadalmPqCgLutU73s59Jr8+b0
1JFYFgj/KbciE2Ju4zdzZuF0FdcYpTns2fQGnytms7n2Wo9z2edU+7FWAxET2Kjl
mi8n3VCNfKp885jYiMj0ArM3t361H2uKs6xnpzB58xsCsaENTfDigKf0gFYRlzTW
9JQUiT3AyvpET2fIlvmAEtcgDrcskT9F9OvkCMOOJekljpQyAK1XQzn/tfvbWh8h
P9sXsfVIaSTBdmiAKgaun1cnlAMKxRdyDOGYw/k6Okbg9DgKphE57slisPVK0Cni
DkB5rSlRDMZixqedUSKxUHJkPtcRsFb1eKA+IyZjFh2bFbkto8K0IPgHpCa51flL
EQvSEs3MXWvYoK6bk4lZWUawvcbsgx9TQ40WIL4qSCWjZhcVlMQt9lkJWFOXtfWP
ia5DBUVqey//jR1pj5zuxs9SG+77AY5TK7m5oOooEHiftbAcdYypkjbIdWHnxLkY
91mFH4mhlOcAVAI/2WJqGAqFRB/cuomGc2D6g2pQv6ROgMzDUYV9bms0e0vK+kuY
yYj54ZNSz0jYz7BaOtx84o2GEZmXD+D0D9K0p6Pf3pRDjS0z194KPwHkvTokbsYJ
DXYTmO/Uvni9cjOeVAstgGiPYZVXIssTeUiWgYSFrf6MRN5MhTt4jXR9BlVFjhgP
GnNJrEld24joy09jkTft7hgs2McJsAwarcWvIGnOjX7DViOM9R1K10IfSvKbajLT
huW1F258XPPbNNq6mxTTU2f08YY60bFqBgcIG14ks/u+sbQi4pCCnu3t7AKtwpd5
n//rcoRMnYjEeQdFdg/Mrw==
`pragma protect end_protected

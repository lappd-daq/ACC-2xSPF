// Copyright (C) 2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std
// ALTERA_TIMESTAMP:Thu Sep 13 06:32:41 PDT 2018
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
ALAsumndcVo033KyBjaBRQ2Tc0Qwj08MKm4TjyCdLkAR87szpHPRcp6A66llNgLJ
xvb16NhI9pz4pFKJasqGhog4BAOEbskGYp+1/2C7+5j80n3IGlx7c3mjWvBta4ZP
c+clLKSotaib6hm6/84EtUdE9bmOa0rIOcVGCKjWsdY=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 1760)
MtornD5XpY21iaa+oPBO83dy4yjBY7bN39WDLjUgGRPzwV5OUBDz/uS11csqo5UX
WMXImwlqwkjf78TGXARpDFF6aVT/v77YjAyF/HTm1aFUY9FcHX+pJVDJEA8oP0YP
pc3wxfcxKcH5xBpvuRs71FYFZGdzqzOQKuv0+1G9etHYLXAwQ7jDILLeDgMRC0WV
DjwjztE4AiI/8vBxNgm3BN6x1vqbDBS5BFn83fCnDi6XGXgCOf6ZlVzL/kmkrw3H
LsKCuODERnfv76USTfRqNEXGPqotm5Ae5oSbUIStyJxYsSdMjxqqQnxcXnVLy/mo
10iZTWcuqI5WQo/S4yqWYGs8whscl/zJnvVpQ/g/w1qUzP8FwLEJAnULE177s9v9
P335cTN2Dw6P8s1lMHAE26Z9c0iorOmeJqjZ5HblX6MaCK2vBLjSiPKvstX4bWAJ
SSB2co86+BWVZMaqoE+ySlkFCm2E6c1ii1X0Zq5gX9vgXmsAL/dggA6/zt7n110C
skYqspoc3z2e30xGPVnZvdy28PdX4AJUWet8xBoJgFPg05CJMaiFCb17iDy+4rCc
4bsuusPTqJ/fg0gTgZVboFhfXYYA8z+U/nd17gfoyd8SY1rpjMT2VMKqhFHFn60h
f9lZPZ2CaHm7SQd/jKprJBDQBD68H65EMnqOHL7PcgcPGYfslW1jwDmkzXhIfI2F
VOp3c5I9zW1Elpii+NXjnAbrSa7XGJLRj0EOb8z1C2EBifm0xjiHd79OVeZyAOAA
2RYdRt3q1iEVsZb5RK/JdiFhKtIVh3NXNCl8WXNi8MDPwg8S78x/jEunle1MlRDw
iOSsjnrJyvH3P9h2jNBKCYOQ0TWaKYZ77s1o9cY2e3T2UrMcPS0wa1I/yfWECOgF
1AS1fS7/tkgjWGBSNfo9TqBOgtg40WEHIGAle3BNzygsWIvmq0i6qoiXDF3CsZUa
zEI7Sz9VJ54A3PI/s2HRYyR1GiC/M5kolHPxC7//M1wXQONfZlI+KLNuGNvmGZZe
JTIvuysRZAyYuJTdq2rlPBPWppN764UShKjIxGuk/8hquF5ABxV5yb12shcB/5hd
7JJIEo6d+ThuUFJ/5Ow9QwLBdn2x6zqICOGZofqsw8veBdg9KuOne1c/yor3iK/I
5FeLP/QM7A0VjIoSPuU6tVmdIgdtaaz5jFXbltCLS/IBwZalYiOov0zgrbxCCyW5
ZgzBKcz39VQEya6ZMPCXa/4Nhh6N7X5Nnuz8wEULjPW4Dt2Q8COjlq2UwKe+xL3r
HkCuNCtp8BQY9Wwkaz9Rg4BaKcQx2hGhathnOJ1q8SCh0xEYHWB7X12ml7upWjHd
yCDL3N4BGDMqPJL67gPZyRJsTYAeI5oMYmCwrDKzQBwkIXJdkejBuZjpzQt14dOT
Hm4rmCEiJ87+hiuNdu3c2ldwqkFRbIdxDs4FBIqehN43eKgwdGZhIwjisZih2Ly8
sUM5wmWJSiosa6to8cwUC1M/x3gwTepvbe8badq+83O72bKafHM/6ZGFDjqTOUJ8
Mg14YsNg15/I5woV3/DT7FSE8efdTykAH0rnAJ8WUiVF6NfeRknQtqWe64di9jcc
iquw9mgievrR/GqkfIW0FqRNZQsGd26wlBXJsFV9dFtQPkRckPpY3yABTr9rRcMl
CfMz9PabnHD/ubupx1Uc/YAAseEeicJYuxblYktaDUpMPR5aiDsLKIz/1Bj0C0A3
Fqjc7Sfmf8ZFZBdlSgMG6etK2uVDLx+guGh6VMC/fEVHWz6uJr5hnAdr9Csx3vzO
9Rut6iz7LdOOSqO+9ZGeUAAyZHH6V/LdZYtILbQxgzCAcCHZKmafPGQxBogmTixt
Tt68ItosfqZBGAYjtr17MvpiX2l43nQ06jvURFyWtaUwjKVJZ6UKIO7jSPIJMMPj
LtyLQ0chOjtQJdwdO+ezuo3mkAU0bgh+L3zS09ToY1wFpmLFO4eBQ7reHLzJ0jRx
H9o2inqYc4pBAcWVnvhMYgQRe26Hj4fD9rHEyy9NvaYZg1lvO3DoQJa3RBcnqE2S
+tGJIhpHX68y/oOeMhuRyAbbTdRnUDDJbPjXaEQ8NRAsKwZWkcKxVF/EW1ZC6mtV
8STcdgOIyrTevb9f/vFEwv+bTt5x/3/ae1OG8Ce5RTg1XttqsELSKE+6myn2Ln0b
jW1MBJqvHc0qauwRKIpbtcXAvPIT7iAxzxY867sRvIKyIca4vUSr0YuX+7oJ8PY0
3qEZaO9Gt8kyqm2BLIiLrsp0ESo6RuPiUAev16I5Yw7krh0PUyXJXIclmkCR3RHL
LDCPsFdCYDdDptmUjbSCRoDfmcfq0OwXw2Ozxhf4vCU=
`pragma protect end_protected

// Copyright (C) 2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std
// ALTERA_TIMESTAMP:Thu Sep 13 06:32:37 PDT 2018
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
g7v+0j79ALa/YOVJstapEIIsqVCtRWONus+Jh5/O6BYBgoNwy3Q5+3A7dOPewrIw
7vlQRXXansa7KXlTyZawK5Yr3X3h6olYvKncaTrxMJELamE1Dqh4wmx/WmxVk0cM
jFeR4sIRmOD8nPMaFdaDaMxh+O0v4Ul8qGv9U0oLikY=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5584)
p4+8L8O7z6qD9j0mxnx1luMgFGsA3ooMBnhNm0HpNuCzkeUujS9ieVLoIgvPOhpi
PmPXLnO2LNgfg1OZhi42QWX2lTinVkwgNPMGgb7LFdD5T2vxD4RwtpEP6Um1z0kW
B6PDub0ROCiQF5aK8UHYa7WEn/4/JkLUFOz0GpzX5LLew1rxH1K1+bGE0EyLvpVJ
/wXcAKdEyo7J4kINq0yGZyiAVKMwqOkN/1sGU7HllYoCdCqDPz848JjQmovmgdov
iU4tYY2YuU+otrh/vA3wU838iYYuDYZRxvS5NTKjpv2UzUdwIPvgIZTrmXasQ6mW
jFnQM6j45y+go83wzltFaxNShOOM8adi5P/xMTg56aNtPVs2XjIQKmb2DNgJPfCP
7l2DOAVNarGgroORMfqIMbrM8BGo5wbeH6aJyGPvZ/bmd4ikhQ9MpWUyKWtBBVtW
CQppEB2LEvYhmDeaOuyF+4h986KVxWwno5lmQpTVQNT0H8d2THxx4n5P2ig9kMTg
6HILnHegCSu1pkWUh0uIwHvwbuYRGLoNI6Hh6QLryJVb1DPRgyEHWld8wQp9oDRD
NKVOT8kpZLawicFvjJpDa9SKLApha3kT5HID0xloCLg5STbYyZF8a+trigp8bf3b
tCVN0Ja1zfYjU+iARIkKA2UQMUcnTw1oqs9OjGmHjwkpU0xs75exlt0ETOzsQ36c
At9Hr7FEkLh68bOVlbkSxGMjaa9zT7GA5VWEIyw8wsSIAecDUNNTMgOJNGequ7tX
gVI+m+67hWKFCzTJUH0DiTEtAKLvfESKNpFqUePxoRfcUH6lV09xbsmSzhlQK7yd
5S8kY+76xHe9LJGHRifoRwTiRYaWIZGziZYGhMIVaotspogVQAxb2ehrndi/qfOK
IVSWmkp85q++ayvuVcSvwtlKmsauPCj4oY0t9s/OZixUFWy7Q31Y2DqC64dhIq32
wPgriqncCnk9iBql43RQWv/QeI5rSTzMLNgLBZJNtWZzuAECRjEZsQrVE7c3ghYI
GNQfLEhZw0bux349nFvjILtFsdr1g/+RzlyUD/CsgIypE4tAuKVfEElqH9xVPsh5
Knw4jHd30QlY2RO6AXZU84c5WJXCVycpkv2mJz5X5kjmxTOd0ri4LdY+VQbcg91u
rDzHgvvQkMlQofNFWpmPe8MDL5pAvHt/eXEYsqLnzAWjCtwdGlDa9ZOrfivROjxB
28kVF9QkmzyIedlEWnbvd5e0W374UerEvqcN0HSlO36RY4FoStfd5R8Ffl3b9nk1
/hAy50fZu545Gc1mB/tNu36XsZP+1Hq7k2W3/EaKNCxLoS6m1mHx3lwedTogH8XT
xdGFE6auXXTaoLe9H6R3ZsKWjvaLOVUhGdC1CN0f7pbkKGR+y8qH5hI0d/7qMCmO
oZCo2XvpH+pL4PBKM2vl4el684zlQ1N1cRpo7mOZ/NUnGx6HUXbf3hrLUAVNHHsx
IY1qouKVzhe6myJHO7U13QLNR/GhSeMQ9z33+ptP8FNKxeAOU1yRXlAjqI50ov4t
rHhU10yxnqyC1vVHtDg5bjJ3Ztdl7Z8TrAzxkZo5HWVNZKHOJSukMVlit+jPJ2Ko
80ZsesB2XQ9TtyOF/8pULcsZg7D7dR55SWeT+4I/vlcK4PgQjsrbbT/LPoREEDtT
TtU2JRg6Bk+djH1VidjZAYcbFELL041jaaiu/u6U3GPFDxeeFwoJNXjnd4aWPRsX
xPavyTkcrgTUo8bD77eNXwMwwCRYBvuufuWJnYMbZLwTglRfi0bDzyIr5PKF8Dlr
JtWSLJV+mWUU1T9gbzj0p2Wg2ysuWoh4V2sz/Ks5SkZt53NbEcZgm2wQfe1hi6VW
vhelsmQNV+paTEB9ZuV4yy4wsbi20DYQKOu2o77ROZuicOC7CS5T2Q+s/Cg/j647
X4dDBJAb7IrPxHxxn3JETbzRjZtMW8X6NxLFxun90/PGzJDgXbM0rYStoH6ZGdTh
RN/HSdHC96lpMra3xr4I+aW3Blben7DPUVngMcsF2JWHwnIawADbYLahrye2OLcx
9Sgt5G4j76E6XW29Xi+qzts5pppB79UCgLKJIQX31P1iAbLhkf8V8RFKMp/aAssN
LqRBqXFL+KpZdBu1pmj9qqlfE4mDfu32RvsnV/gvADaY5OLmJUf9QaFMftPtEc7c
pNfJSLCC4aM/jMCFUVlJZJTBcS8JRG5kU2LuHtlLV5BkWZ019fOpM7jjRLdgCVm7
IVkHKviwFQha2f9sdoAIqU4ZHKGseVLAXKvYZsiylgjAW09AR+yvHYE4y8J6jXb9
MwKWl3ztFvcHUzkGLUWV4DzLIdNEFXd3GmTtowegp/byuz423wXK9mVuliWx8u8V
jiuxAFBsvMGoZHhmesXMt4dJKH9WzktOkKfL9yJ5ssSia+NKamQ0RRup9/fPrOz0
WRZV7bHujXdkvtUGq0dAvVq5BjOH2o1HeFnK9M4AR/VQQXipDoXabc80XkxThGCS
UUiKX6NugWp/MRGfNpme6b07M5DJJIlkMjJw06AdKRBYABv3yyG0NEoi7Z/ORImS
rHPHpLHcMxUX1bnIJYqKO/B/f/Rb80+MMG49ndPY2EipSkREeBpjMO6BtNaRblCe
GMYZ+QhYG4COltuJq31OMl9dJV6JFwnPql/L079fp4jD3FqkD4K0o9iaFxixVtsI
847w1xfSs2tEUwEhT6VuVLg2fru9KcKaW4xrpcwYGCuZISxMYEsUFm5e1h49Uxc8
zINIcHi+JQLgu7+qAOYWLVIqqbae3ztF8Wjodup4Uk8iMdn44TDlkHm8q4bO0uH+
Z1ZcsQVY++ej4Igpj6tVbT+lOp5icNGXlN8eh9u1n8C5boGA/LKkDRz9Km1gzHiH
teF+podktKE1eEGCmgHWfMeZpGPuhwrjgz3wZsbXsy2gdMHAZcWB7SiA1/NGojsY
6IjneviVruUQYgMoXLEyBU6FgF8e8RjRYhEsrYqpdX0xqOqwD6wzbsnl8ytbuKYF
YSVsLzh5d4MWQFO163M1NscsJnGYlO0rIkFNhWorpVehnvwLEyKApfooTJr6v4Zg
cZDB/H3SvrJP6/YDECMEnMATSlgbXSDjMwXQWgT5aQXsOeEPznJ6MpcTR5Ac4/gw
/vztxabEsg+M+1j/C6SIfOn+BnH1mYvSt2LJaVrKY2JC+hiECGWiLjaq25Lm+HOL
k9UvsWrKaOadHARflhUOmlGWM+FK8Yw7NKPwLf5tg34c8uIC8FAsVHKU2hLqNuVB
ERhIhCyd2WisA9rtPclj5Cb9Aed8I/IjD0/964T+DykaueTum2h14Xoa7+ac7/sR
47kOEjsdrh9zUXVXjFlFlLHoB1FYcssOjdBDoRNyOLYay/W96ZMBZ7eNXYxGDNsR
ZOduepa+Z03EGI0B7eJHYb1ADLUF2vcEuRKA92HI8v4t3SYmLJpkK0Atx0CDMbs0
JFV91UnJNl8bzrVrNhxMV8RtOz2gplTg1ZKYpUU3ixWgmREFj2onFTagLKkPnULw
W2FwOWSv+2OafcGnCvfmpPv9ODbQGlLju/GR2UKjWVaTLONxDNysXN/b+PSIS/wj
dCqNYddUJvlryATYvfLYtFb4VjrhfRCFyguvY2w8u7bF3ZS4SQh42vsC4/7C/r3G
OKKgYnzYuXhwH+5YT2CEOj8vqIiO9ipzaq5t6enWbAxHiIInHBr6crOcWwmNZbOS
Y0Q9Xo45K8KG1LnnVCXdzV5mHQWR+cdzlOEk1IsEhwZUT9EGo18wj47MNPs0ztfJ
dnF/4npxB63giY7KUGGu+ailSHGGkyrmYanUpJM38NpUpVnjIvTqiYJlmHNgyCPf
saB+WbApDrtu+39Cy23n0xSGmsmBKwFGUepCw1ou/BmhfET9TBcZ8Q+SQGzdEt1j
nouDqWr1hV5hjkQ/R5HaaQyHMfqvjmi1xMy2CYTVROXB1Bky/VE6V2NgAO7nOAMF
lzsBFuS9LzA89fDWIJ8iXb1SSOgfb5yucjN6X56eTLMf+PyUU7aqbPTAHD3icUB6
/OjkrNihkuK67oy55cHyL51I8kw+FOmlFQkfCF0GJWkS8JIUEfLnpUUFkR6TLKjL
PEcNf9NjWb09Tk3sGJemEVt6rYZaYeb1Y0NX1Rh0HPG2Yu8WqK0T9OGGG3ETkUmc
6HKzsnl/4Vc7m1vdSaD2+dGs20fpa1ZrrYQXYThPLtnRLacS9cpaNbBQ+l1gq9UI
y2E3rkX5cH2vP+NSiLLVYb6LzP4aPaHefDPW0KH8nP5zQYv+XJ1jsdrL7I7UvdXF
bV9Bh9JSc7xLmL+qmGga+8tS4OUhfL+YFMiugn4SufJU7rPQkba1WlkGKfHl9eHC
p5vRso2L5ICiflO6/hycRbbfw3S5cxDgEA8CaYucn8piqcHqQbiYZpM96uXAv8wz
cFPZqHfCtrtMs0KgMQB8wGFyMGuRItMerBHQBJM7KgqnOFiwWY1jYg9uU4+spbFi
v2xQ5fqVCtzLTQY689mIlT0lhhUF/Mv7EWMy23ezAxwOCHM4bKXPDNF7eJCZvOSY
yYHLtZcYf0Jl0JbOOKynGLEeVZCzkOp8CWWl+5EPDDPi1K5nDkrioTrkRRHRMxBC
CwcTaBSE5Dh57NIJXOpJDu196x+rI+KtNKDuF45u6d5aNPD8rpB6sHnzz8xWsXr+
kQQH2CdVk46phWWu2ThPZDo3zqDr70XescYb9WPudRgRpScGkK2zUL58XZqoJnV9
WGzbyzLRyri9UVrOzMaLoK26Wgoznof4one3HKpjEKglkJtIfrwg+1QSTcHb+qrZ
eixSbIlOjmKTDE1Izt/wfLQmxfiW3oZDxUsgVe6J1b1MWCQm8xS108uiMIuy/sfA
RoqImrUpjx0jmzUCHo6cmTZ2LjFSBLrfVAOVauMMAvhUT9RwEJwuI/DzSPbIJx1g
AGk+NhlBcHi9vNcdksYF+FK+EKfzV8Mfzm4UBF2s/HRcihpfzZyA9IIP7MHa4dK7
jGyP886hdLDWMkBscwyKKHy+QEU0lB37vq9O1aWeCFh3mODustVSYizPZF9DYEDw
dA/+CBEghQU8itFPwz6nSBfzRV87b7n+ZWdFHgf6grfJDST6ZOGR9ABW+h1LrHgT
46/mnkQUwYGujprH0JdUZQHt0Q+FXELRaqm1pefBS3/F7lpHWcmX6PmwZJQI8+R0
czWiFHGd2PjXEJTOkxthazh9lC3O+c3a/HyVtBgXODb76QBVKEZI5mon15WOraN0
+9X15wTXsG5vRc0BtSPUt1m2QvruFCl3irvnI8XIkXHh/mI9Hq0odSbFF5H/Kxne
4WuaVBKHUWs0UXNOhhq0VPqztBvpmrXhYwLQQg8FzQpgJLDLAYcetZfCl3DdPTtb
ddS1Mtod6tnIl/b+f9cNrGC0m8GpVcS+CfxdtaVS9vp6/lNqPUDOgoWoQQbwBG1i
bxMIdeVanxcYZEwg+Py8jHAUr5yGltLMjpthDfw0FyTp+tBDmhhrod4KKaX36jaB
v1JpKLO9EG+uwhjYuCnwEjfWf9HmGMQcuL6llfu40sN5rEYiUunAsr1tRNAZSSlx
C0vpqKGPh3mRTVIxZL/W/1DvRoaGY3NwVymvL+zHDEbxSxl0Vo7xmCTBblgzOEfB
6mPzyLtVPUahKwhST03CygBrHqga59gOCtridgIZ1V6QtAv1BM9xwn2KL4PaCxKB
wHrh3mJ+fWYJLkXhcqvFEoaDp0TPAYEbeSIan00zbZ3TvJk5jd274n89jjt+Xm5t
9LbOVsGqk4jyrFesSYcY70a/Sw2FxuVTLyYa9y2LQwL0bZqfxPX/i8eLb3C+VXUV
baj8+9XdbLdyqZm3ES6vVmjwnHWgcJWz7rBKdJSpfRQQHEDsaAiYei3L/81lHXDP
JmrC0kug47E9ek2tgjaH4A7LUChNatGQVaFby28xxnuZAwAZSuPCUgBCOldak+Xe
Y1VxWwYTQkd4cRRsTASnMyHBQtf1AMCulOqi0gr2+Wo4e9a01oDMOBmiN5buxZSj
o7c/TmJwSjFgVAET4z9rjDmikfYnIBeSVcXAd+LuOpqnCMnZZ7BNl+Bdqtzrvrbq
QS46hppv1xQ7LG/YGcbUk8pxwZrd+sEWJRDwzGB2PO6/OdLCsibQWPht1s1K/Cu5
Q6GjWkUbY+nMKUtfwxyWH8AIrNm+rDYsdlHvDPulYsmqMFUQ3tQOaZ15gaHbNhXA
5Tbjjq5YZ/ssjPvuwdRCgTajRf/OBmAN5CSaFemXC/QY/yMQ3//gle6KfrV7DwNP
M4f7pUofkwX8uu2Yi30Wnad7pJlF4PXZSgcB6Mc3f2DVSWEZc8TTC577JwXk5qv9
ozsnZsCf6kxvXhxF6LMc9keuNnu39UBH69NtMA7OewDsno4d+gsvHjh7lyxAlaLj
PB5a1WcTp1P2b+A4tdi8onUz6/60pGyWD3YVpRITLRWAI1EL9PIEJNXVHJK/mI79
sn8yWebrJrR5nEI1YggLkizLu6M6FmydTW88fWhnr+gSYd75flHRZVFB7hc3MWUn
lrU7KFL+QbHB+KBPPA06H7a+aBhlUo2rMTP9fwfoS859fY7B4Qxba2Dfp7FgsRby
zhNLDlbHXIX3uj+bwPxmGTX7qEXFaHQ868XqNb++o6AroDhjuUc5g8T4AKQVMJx2
JS1kecMEZ8NQL+sT2KX22xeGy0nn9sECQdSibAr3p9PPAoxwLlYAJ4jqX/4S1wd4
8Ofoe/wOVUbKguATTpVQmr/8B2sxfSsgInrknicwEw92ePJQ+TQS+nAnGzUH9bVX
ZV0BGCatNN5imbaX6WzthXgfMUrf4RSSkRqxaiXvV3lue6a0sTEgq+nu6YoQKCMw
SlhCkIUjTP4BjuRQC/zBb+0TK7tOUD+vwwJneaEhQ8l8+6DcclFCN+XxRIgilHR1
SIs4/ZfWHyk8dGVrftNWb8JRC1ZeU+6AL27KxCZHi4onJkpDigntJ4nMzplWHcPx
nBJKv/Nn351ICwBjEqPNfWbNas2Wiuiyn9cwr7lqL4dCyHaBn1mOHbgOnBmeGjL/
r5VXc+fGz+2x7XLb3FlGJC+MqiloIXWPumcbyD1ZQ0hv+y54PQwzFYqSifdyLJd+
u9SHhka4GCMnXFJdLG02dot9lId3jlr7TXtwJqt/myXapBKh/qjkncg7XSOv/vM1
sxLcIf1GM8I+VCCwb+C6zp89UfvfLWiEy9U5vee+eMG3gUOoe0IjW39y+I+z4BvD
dO4qu7mi9QegYlxZ7XlZKj+NFiegSgBx7J2SEa3WfNZJZf/O5JjIXZWn/qKjsufp
X2lQAvCB3Nf3QvTvs9LeT4WznJ5UKz9ZcCLrTSRXISqWUtUyjoKyDD2qQbCC+Mko
HUxHSWPzzzhWeEkmFdSnf7szfb33zuUrxk7vJpq/UrT1QV/s9f1QilszK3f9+A1H
npbGUZ9qw7XpOxGzbPPeew==
`pragma protect end_protected

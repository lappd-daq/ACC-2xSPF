// Copyright (C) 2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std
// ALTERA_TIMESTAMP:Thu Sep 13 06:36:53 PDT 2018
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
EdBRBlvThLt1VYUd/KlTqP670UqVjbOtAiNv6tYEniBXSxQOypKynb/2Z2AtPq4x
8p18TQFdxIxBAYEKtb8LMVexRfrBQ9x/2xVscDXkeAp63EfmPG8rHuLI64V9FxEM
g4Tmi8p70VJQL8mvO4QsQnVUJYxwxDtNkivkp8IRa8k=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 3584)
iI+py//5JKOkLCBonVH01C9ng2LLUeczZN6parOFtUwSjC0wxpvT5t7UFXbXqi3j
Y75YN0wwHzudRx3q+lfzLsKMQPmzYDSuNVJuCF533evoewhryHa4kpKswTolkqwy
z3nXhMGFAhSlUbWrVRKOT5KbkkPlIcOAqIkjdZR/fnCUX5jBqcp326rDLn1Jduq3
fxThoATsl2Fz+D2a1vNk3nh1LtyOrbfDdE3V9v85XzKmjb1SWBtuAbe/fHtJ0y80
z8W0rN4yy9PRhFjQKbZwcTyDMFqLEuiI76Jh7p9230KLwLzVB9MNDa6OKB74mle8
R+r6MD6J+TDDvXyNpgr896/J8hbnC/oARf68qIsul2B5z7Y99xhsQbqyt+UyDwQp
FgwTeLt0toj74K1HIIW3KYIEJ/1AeyyfDM4HURT7T99v10x47c8wRGo3Ory+iy90
FNd1hF+/v9O8CIN8HFaKjoIAHOPSyqbhf6FpJ4V3EdCNHcEl2wqgqB8xRx0qA6o8
gx32PeK/sAePNx8hhf94Kkj0d77cjAbjEy2ebYotwGOQJj1FSt6nhgGYV2Z5k16/
i7m7B/xl2rGSWoZrFNiHxczbztxw/uq1vhc1V3xYiN1XIORS9fbZJvgOo+Gofgk+
DaSwfeBtqXeEcAFqXwRh/9zBMvdt5Ysr+xzh3l/pSwe0lB41faiYu6pX6vMyYbhj
Je/dyBysecepf10gfVitV/jfhlUJ8S+ul61kEPf2d2ipsgjH/NEDGsMQ/+Y1sEe5
Sp1xaY8qJ6BTQnDmQMOPmKUtiQoMGt/OSR4b1jDQHkAqZ6uV1c83vqzDaJvkRDTQ
UfchsdCg+rafNfvDkEqTePFFaBkglVn+zRpYp+FecC6wKbxqAmK7UtKkHnUKgdOH
kLzxR6vqDZo17bp0NUj/e0mnRamN6Kjy6WGjwdDEP6eLXthoEsOAsqsFp53Z9HxH
FC9nbw8ZrhPUw1WKzf27NEe4weWyRqNR/cYt03yzh1fINBQYQ4K3XNH+BXkMbZNG
Go/aApqx8KsIsti5wnVxAz99RS5ZPVnLWkVwqxorkhCRtojgkoAlYnPKRZdx/S5i
wsPB3KsykFJkm1WyqgSKynBKM9wO/EZfUmmKib3dUQX+hjkP90fi4XJ1ZyKls1Yn
0HxQe72mjKRBTUIxp9uGLqKDKqRj8+my+/EMumeoCs+oPEu/6rMKdm7cqK/USsoY
r0smFugM373mtj7nljUNwY8c9kM6fMaEUlcI40dj6uK79FE5MUFA37sMRB6jtx/P
+SamY/JLoLUNGpzYk0bpqnVUBSdVmcsmGBN9Ob7wtZ9X3pzsf/15dbi+DzLy/fU5
XpPrUktrQ84NfWfVjFAMKFPwU410C3uHdS5H/pL1GrBUF9cxhp4XqsqIcnfCbU5B
UFEOE/QYruoWzUI4gxZgz7+UoMulT60R0RzsGMfCcFe5XKTmhkOdeU+aRKyzb/2w
SPShGisazxl1fmLK1l9mtOpFCrbakFIwIQroSFSVk0/loncvsCHkdqU7400iPKTQ
/nFSXe0Lrs9a6kBdb3DqYNdELRMr/ngCAGJfY2ZZeKqZXrCOYuFmAGvOkHmPOKXX
DRScm4xWVR5cMYApqpQhCps8UdotyRBCeWtRf4H6O196AWvaskFlZWeaPdih0m/m
jYUhrCPG8gbApmn6wFfxo36d0AC1IIi/7UFXb0e1uONJiYjLPIVHKbN3i8syzRki
9mK40qKfPLnT5LbzuosEbSB8fjOlO5W8ZMkXF4ZOw2M/lheIAf0dyNNNUbBEq7qu
TsZCFAvW4mXfP2SPh9RLyNGtOPWkq2KC/H/ncGJa93W7GwIo4E4DOtS4x+cFzf/Z
gljbWxNDji8OtCrRy86qxs6KwuPrkrA99VgQNbI4gAwtQKHT8mhaR0RuSO50PrNo
t1myCovsL6ENN6LyUznMss++Tf0rk8+k/+BSWExni3MO//hlcXGuNRLXDFqXDeXu
ncGhmCR0m0BBctD4tyhy8HIMVbQMIKl7x+kJxKxMU7Op3E7zsYgZb1lN6rzN9ZAF
kjgHP4jqYxpTwThvztph2s1/yfiALdazxUwu0C/mSh0lqinZKTzp5GVfcbrf2APc
TTIMqVOrPkcLYDcuYez5qZQXQ+FwzlmbT0qURIqS5Qw/h/CtdQSvl3tdUgrAqm1p
FsJaCFjrKRahZi0CNyquhrE5gwN3v4nDYEu7IHvKY8GDiL9f9hyOSd1MbGryKJ8z
87zlliH+eR4R+klQp+dTczWLlSGrSVhedOw3g7hxk5aAGs0uialnPn8Zq9zCkSae
5K9gNuSzSG+xhmK3Z7WRa4pmn5LpXhp2MoLw8Ao7wh942rAcx0CA8aU2FrFD3q6G
vlSbIK9J6l+CyAdsD5j2iEQCqIIBayS8iV72llBMw03NBYz62LQZ7nI+L8+8gp9C
2Afo3LJpSUmTMOudnonADcciuuNyWL7iYeIssdDPTVptWdh7ybnh2uKEYt1R0lqX
Nb9VJgSaIMOFkhkIUWqTIsXbBCuZM/ZO7e7TWTMiWCZcIpA9NuTwFptjQjatSohu
k7mnwoMa5jZlwQkwt/fhaq9/+7q8oAHN32XygHpdlnZnDgXB8myHHrWK8sZ269Wh
LN7iwpGsfZkG4xkRyvATgJthc2FQeUUEzmG7OZKL/+JBwG74utapsr+AUriUwxTB
lLu5H73b946So0/pPFq15krYpVDO0zHdUqFE9yE3ePjoL4KD4GXgrqpggR7gsPYj
TlHJnZTjRN2EOkxNhFD8kzS2+jvOu6vmZnXxsTM/iCPuC75v6chEs/iw+7JesWWq
cEN48BdsvhVTVFg5U7C4v0rtn0QAnRsUPU33wL/avk/LWPqgVlb32qOZnm3FHgOf
WdE0DhvoGMbTnfOD4dSCD4FcHmZcVGzxuQJXdBWOYLRVUCwqaklehotPeWSsd7RK
7EI9twqqNWDl0NRt5IJ8trKw2y0ruIASiirDcXXqssGaeHQy1His9HAHoujHPwOl
+iXm38Fq8UC1nPnxR4fCDTj8MPUUW22p7zt/2FjGIunl+m7TtbeFmy7x7SYiWGTx
eYB/YPpRGNzVMDCOeac0ZglwM+z9CTsWXhutE3iaooCcOanmdoBy6oPAYN9dHqo1
7KaNq+/+zrZiayIlp5JVhrpwmdqWJgi4NuCLffLgdjEwpegoqbHikD3cfnUDdhVG
eUaS7g4eTeEZZ3bX6ZmxpZ7jVPQq1PjRLUQg7CEkEO0+IQd7aULWOQSNi0x13Hz4
69p/N5Y4dz6a3XuppHmyAas5vb7JQd/OY5s7jUNSqxMSTToscycZVCDC0GZjc0Ib
8KgjHwcofU8lB6f2pKLU2np8IzY989w1oP29dVROBP6UMuTj+brtbqyaLrIRvDff
e1nFiQopLtTdghvG+dd7HriRfJS8xdI4xkyvFziOj4ChvX3/GyGjxsRvoW0e5IJD
rw3/ScU8pTSR0Eg/MCkzF6FZnP+qRbO6kBHMACsl2pj6y5ERjbk4akSXlnl6Optc
BoTrwN9O8XoPsCJo+Q5RY7BJLmaWWOAC11HQ9qpePgUe8obIsOSVVB328xE6y8Al
f7A0iBg0f4qmXf8vuT+BO/g7emdgSfKphy8+rUILNTYp4/1TsqDiSw7xlAFv92Mx
RSdCQwxPymqw4TH0suF/hsU7rc5s5PmaRtiZzPO+eTp6QiIx2LMu5qAuPQyzg036
jkGa+oZlLW9BbvipnPsfmmvut7yRN6XYlmkgfHcTqoW0NRCVR0hfgpT4cNCHUJcf
arJMe86sgCTM+oEQV6GRPUVtJcUpsfQL45dvYBSbnj5teOnvP1oCTdwSvK4yXT8U
w4JJtZJGaACL6/DwYzBYzxRohOqsUtxBagVzdnNcPrdDMU5G9tI5NP2CkDam4tTp
d90DhwRsL8oLsed/4cRgu0NWt4QMDKbLsRKzaHbF0JgHSUarUNAg9V50VgI0ATFH
tE04JMashtBwS8JP3U6NkGdIJdyv4bkc8dU7hhogPLllowJ+xWqCWLVeHS2ymsm2
lN9BxEQheP0SOieCmpp6gEk4BRn5QzDKyfPY3Iir9NOmVGDE5tzhpHjoksiU5W3l
BOoWnRmMCHcYhL34u7cP44aLTIX4gRJVaXaQEBPZcE0e3V4y1b+bMAyWz6xWybtU
rf/svPmLFKQ05zm67aLyBilxoqURN/ouKz4SiKggq669Y0sKW+OHnRyGVVpEDrXs
pG6GPkZ6/l0BzhNyZAUNmh1jM315E0aMMoprmIad0soZABgpUq6qxufuGv9Xai8F
RuiiKMrpha/1ReOg28Q2RBeHH73g+9cEuv6jjZltnd2uN43cZMVi9WadBe1hsgmD
CH6NwD6FA+MAA3ijJwNx1GRQOKZoPSj+5CGk9OVFB3pcw6nbqBVhapIMJWyK1PQ9
wyf9w0VdtvHoXNVLwHx1CG/eiZct4JYZwLRq89fpMw6QSsAs0SRsLIp18LfEFbbO
W77ZzLxeHtjnP3NSstEU9QlsXF+NRljT/pB42JfmcbvrpYXE6ADScQ3KmwlYLMCa
3LiotEq5EySY10PTMVwNUkeCQ2tUJMNSxPrueTAI89lGKKN4mX4QM0Zsa8wRsiZp
ewNNPI8lnRHp0jLVkJg19aPUoKwH2zZapYB8aSd1/WnbBD6WID0rJENKpqKCYAKu
PqG0GUU0y00D3zuJxMjXSWO4/zF5cKYW4AvoSMl+6sh3O1MGgrH+DUJlhiyN/GOt
MNNWohOlpiLUweRQ8jHBwpJiNqDGpg8y+4MyK4gQtvA=
`pragma protect end_protected

// Copyright (C) 2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std
// ALTERA_TIMESTAMP:Thu Sep 13 06:36:49 PDT 2018
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
QMCNXCjmbiTX9Kb/ZE+SVVeQZTZ/fIh+NJkeIOyZ7Y/QaAwDDguYCYA1l3btHdlf
LJ/HDivxXN0oJs/MpGtPD+EmHe5nUJse2j5QqK/DooR0yiM5GCmMitIW+oGKmba0
0P8c8tbr3gxoZLOM7DZKEZP3npBkqXFlobpEKpWotTI=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 17280)
9On1FrVPWp46d4hxUGsIC0uaiEBprYrRtVHgGPVw4ZufaA7WU6J1H/HQ8J2mD3ze
jBrbx3z0SiHu3hAuZQeP+9edOfOZul/boSTxtR8anZGlpMAcGXEzpxYwvi+zFWs0
sul+TXDGiWblIluGv5RfYSq/c8EQixTyJIXU9VxrC3Boe1OPQU70AIvnmMsTcjcV
fYprx//tXKFKuW/WVrkL0CvZEjCfkqigp/DsfmDt7Ir4J1MiH/79harGSSjsxIzP
CljMWB7CjyAHUbEzh3kEiJxWHMzm8Zgqs+a+gwHOoSZRLUpj5o/L/snmjl3gYpqF
czJ5lGlUh7WxTAYXx2vsN6+LQshEfL5qquDS7ngk7BxYP2BE2b1IDe7lI9Ge3sWK
VTcRneD3OkG74qTvkeU4RK+UGgYkvQqOftW+0W3q/fo6UzjvKaLa3+MinXqaxFXh
Rn+OA5nt3igMcMPotvqHQdkEWndOOKKqxjHD6JtF/he/Vt+3x7yiXdwtSYwVd4Ri
4nFs1/497bSWurWZpAJPb8FGsLIpi8eDfdKcF7dmfjXp+7B6Awki66r1XEkYVHuZ
yTBgtsog1O9c9x+B27Pv1bC1ZolDjkkN6P9igxlsB42711KD4iNWWfo7DrcOqqF2
dGzFvqLd9OThAERsH7ZBRsNWtwgpPqphs2D0GfI6lCaNKW0u64ukxkZcuxAM5M3A
Z1o8Uo8o2hVhUQ5UAahfG+leyTZ9bxE6uW9DTdRbPdGPzWSHVeBf2b5MwPCqOeCe
6bJasS4OO7jnG0tTuVaCJxSUFBcfKWz3XuQ7RTJMkKTUmTT3QHJZKI01xW+fKfj7
CtLFugWalvYFAutDLfJY5Tx7bcEXpmYBicg/QVlPHYRREx/MVNIG+Y4gPiNZmBoL
cZTuaL9Tj4bKz+92ru+0KACS0xxv14Djvn1m9AxZrqpgeVBH0dRzj3/xnhbNQZ1V
cAPEAf1BCKT1aqoYZiSor77fV/Kcn09Pw6dvtOeOLtbe9NQny/IBCh+u3TKnD5jg
aO+/RyKM1uJaMFFgnBiYsrZivpPjmjXQiuMn6gPZqdZI7Qen7MGDbMDjb2emBWw1
W+vz5IaMlZefIj4fVUO3TIv+Ohn0AgjGFhI8H/LrY/ZM5lafqYDa4+z7NvHWw+P7
q9H6+5zOWTJ+LrUD7OfMmccm9oNiT8AHU5xgBbGSx4THybs3T6PDyEVpjkEaxeDN
pr7O7esdzMAjI/k1W9PQ6rExKN3JbGlvZP4RJkbUVX1upVGQxgdCCWmyZ2ThSPuE
XVXwjPxdDyHx4RduVACfJhyH6qPrYFEorvfuVATdGb6aB1wf/u3I4YKIfOaSwXLL
277aF/tzHLkQcofH44kjCH2cP6VXDvlHglcFinH5uO83Uu07/Edt9LGWy+f41IzQ
TwBViBvj2k3xaQ4rpYjzwps5mrBXuVZPKOGPTxWVZM/05BKqFjzoiI+X2Z6eqjNn
E1U2k4rxyl2bCmcnKBdkXE5NhJperpv8ed/feJ1fyoF7UoLHNIp67IsjJsaEsMIj
xAbcPx0eYQoqKSt0DJw9eBE3tt6PziGFHkBoHxLpuoIpvHBCJl7GJR16ex2AvM7T
LWDt1SkANpvje/W2+cT5pwUTgv4Oe4wwCsz8+tRBSakjn0x9F8KE0XSAHdwBqLkr
izKNdNVrfBlcy/+UwXe9gxt9NN0XfEl2HJ5WDMOUhcRmJ61J1iHgEHm2oQ6UxGSo
A1S2r3blxfoKc/cLEGrcnGiLsTnsKqbt3jXtBxARwPt5XBuXtVBLzT28tkj4y7X8
nCD2Zet04CpfY18mgvknlc/OJZXevsDEc6g454K+1ha/DYIOaQ6dUjXdLEVOEzgC
UAPnlqNcKZYUZ0o/u8gFljf2XQ2PKdWxrnJka/pdQMBtLH+HPPUPbyhn/dxbUjEX
IUrc9SMW7eb6fnuvo2pyaHloKPEgxUaviUUwaD3OV8kgDhdR9m3fUyvnBC7AxAAM
PvedXgwmdFFawnRw7uBqNP1UK/WnElbKuoRqvr+0vchvtJFtbv5vGTt2fBb99F79
77nEo+AswiToV5omjZj3uqz1nXBsTXEBmJIbCZY45bcOBGRsgZCiZpHvhhH/Y6oQ
C7J1YHB1K/RWmfaW83BNAqlqWPzt0HyukP5x9TX9wjoGIO2C02pwV75naQUvDAyS
s5C7d94e/DTBekQXRWOhcYiq3HSXuORs9C8oQmv9btFRmKErEXfsG33AaP9fQbqd
OpLZJ1VR/RvY657blmQNL0itIQYqxR+wX35D7view1Agu+7P+nPVPxFJ63czRvQy
UrOz07kSf7HT/NK2zTnfy0J//QAfbotljGZVQz2q9C/IhShU8CyTGufuK3YXs895
loqWtkSN/GcrTAmzJ50BRY/FIxdFiWe4Ws1VopYktd0GVqkAdWzwhFVMCefMGm8i
G5oSRk8XuQPe0xrf7/xamrNv7s4uXex7dZpXpdbfpNSUkijLJTw2cUeimNraFvdr
4Xxq38n9h/cPiidCB69ZmZDabAvQlMx+TS3Ha2upf64ltVjzplakRo6Cf64koDUF
3eQvTWrpajPnIE5m40rCF+CGtBgALnJIJNlZ+ucIIeSFyYdwt7NnA3+Vq1ARgehU
/SRPB8BsKTh/Q8AYVdoBhh0KG/mUOZ5LgG5YUUoU/CuxCft22F8YgyfpXrZGo2Is
PDKQcgKv2sQnLWJdnXDbmzsbguhLb5N0NxgvwC5TkojTvPwg3kgZI8qa6RsTWMBL
83aardwJ7v14FELKXyDSL40UQHBJO+xHRi/U59HPyfNwAfb7ahrwK0qDgWP/azEL
WdRwg59MbLiPj4S0e9egKkJgZdA7R8IIxuiQoMw2NdqQUXnRJgkQB5OuSX3bJqqO
IMg4RnMNxt1zv+LV6f+/XpJ9jABf3P8xvCZNl0sU8kPRudbXmigwUyrf5r/Xlf7Z
GcW4daC3GrdKrPw//KlzVlGaCpGLuF+01MX/ZHH2Hz+rxVnvVKRUGK2ngldSDm9i
Eyh2yBDR47sYbtsuVEKG4jEtRK4MAYGPHdcWcI9yj9EFm+AEx0ZxbM9vMYzlHAc9
+porzhWKDa/DNYeCfx6U5KIlQsazmcoNjJBW7x7iO3JW4FN0L5LuYZg4fXvaREn2
ej3dXI2I1cjqzCLy2Cvg+5IM/P0EV4iR6Y+CuegShw/HVf60fnZooNXwUCEyDAe1
zdSU5MfNrr4dj8/b8l7LGrO5CUptqeFa7zb/ICOE6SSlCBj9YPLWh0EMTKxCjqhk
pm9sYIXh3O02foqmw+yzWCxZW54SZ29wQ1T+EF+hvZ7Gjo4m6MRCtatUwTz2SH34
Go9IoqCArQuf8yWCXnlCXhvQ2vg1h5OO2YeXh8OLc1oTZf3NGX1TQbBYeE+4mIng
LX+nHpIC4ZrcpD00abhdKsUCurOSRH3Dm1W8mPl/si3+78ldTMopAGzkcBLjV3jf
paHhTYNW57seKJ0kRb7HaLGOfwe62IZZBE0d5xyvFiWlyA0zG5AxYjkAWV6P4VY/
XLL6fCcm8sQSLlZjwKPvg+tEzQc1qfTfLIxff98BvVp/z7AUedkxq1mFMTfXoQQR
3j1JQIYIPGh3PGxS0n3LWmgPvoEThogj9wVhXQwZ+vYHrdC47MMPMAmCq1u+KV/+
B37dMG6SZdzdld03TcneO8lymwqdaMafhsXLjwA3tMyEZblRtwS+xsp2JdIME2G6
2z5TcPQumlTi3Go/TzZSgVWzkW7WGwYotF4rgly+/eSh+cWNwV3SJJY2IsHql5x6
v1CmAR1fcSoRXNX050RboiMSQfvHXgheEQuAzbqQ3ly1Y8nM/lcVahfDpUnVYdQs
Z5nSUua+7ezYoWKGAmsgoExCx0taUKR46c0clpcu5waT1E/EYCdymR1m0wkeykV2
2u2icOAsKXyr0brCclz0QTil/9I2SXZzl+xK2rPDmoZpUsaNKZZ/RmOPWnsQk/Dg
COxOc2pL32gKK84ch9kN6DWH3PdQ5tU6Dgby1pNYYaU1KlsF5wSnKUdQ5Ix1WlZt
v6tqbJgVwdTSuPepz8J4kDJ34npZFrQoHssNk9aC4Q5hp4+3mm2zpFT5ytjavhLp
hUA/nai7qdvaWDbfPFDZrK8nRXcMB7eN8hogVEGfmMZBCoo0CdksZH5ZrAFrxCQe
SeYrbHP27/rv5BYkg0mKkyeBtpfQgnqkZDmObEqx5ayOpwVDqIfafeKIYg5GKL9A
Llh5r5HPIrsvdF7/81E0cPeKD5MzqlKYVAMoXQJcq4lvbLNpq2E9bZQ66GmyFbV2
ZTH2W7O7NLzsmd4tw7WCMOA0x+8hGQHWmWRfBuY4TuRrkByO44e/qVmOSGNSoCzL
E0+e5dm2t5OzYxs4gDqdwIrP2+Ui2oBjSxeL8z0hhzNCYvfcNIfL/TugwaJnN32V
CxpztmnmEOtSgqfqZyLzaXVfyVHwndKPoJx5wJqpzsZtu7MMwWqy56foorSliAAU
W95WKHOXp8tAl66Z0nu34NDwqiCb/ZBd0NO1e+BWyM8apzHbx4sD83rKXcvPZyas
dv+4HhXm9oVpPR8VfdLkFgiGzBXumVOvnCci+3RKat292tF56ox2kjwH7/8Nv1iY
IzBgZYCOAnJ8+h1DhSMZ5MhmLr46z5T4Oa2TNVSiLaaDbZBtlUoC8LsR3ycfsC4V
6jnVD+OFuPzj/a93Qrp/MBC1jryOToluXvbxicyUWxL//LwupWLUxgYLY2asK6t+
6cnpt4af4X1WIILd8bpa17eBd1zknjsBVntJgykCA35sYCeSque4N2YKR2fQvotB
fetE6dKHiidi8+UJoIU61YCUNxoQGjdXwI2nVh1ozMH/lbP4JPvNq3GMV8Xyok38
TXwsqFDMpVs1ZocWH3b4gk0U8aLTJURp+VyDkuZUJWM4HVweHzHYtisdZgF0+0ZM
VQWxGPL5J1Pfk3F/iWknDg+MW+CNUCnT6GLFpTMBg/d1R4PT0QxZVQiwbbJjOtLN
1H3jVFPWsv+KKlJYY5ADKmOZUa2IONgiDdPHdAqIi020uTjbw3xdxHlerxUuSkTj
wpMj9xuV1StUqNGuS1pvpLIfU6+o0kR/3y2NKM9IEcyyXi9h8qGSi6FUGZgjZw9S
fDdUHP+jKOpD+E4n4ogp+TWjpYrVP4EmY9sT9s0ck8YMeqEAm965eQygr7GJvQjT
w9yEa7k45Ufd25hcW+QudO2XzlVPLa8hNA1XdO8e7XkgL8lqDSADAnzqiT7J61iO
MKWz3M3dSV6DfdZ6ajFgY+ZxpfacHSgfaVfIBXAa/qV5Kj4rsWJH0ZFJwH514RD0
ttCYgMh+ux7IXZCXN4U5Ia7uNlihTRlFVM761m775FZB9Tk4BIjWlEID214NyPaN
bjduHMxFqHhfZcsgGLCXG3mj/ggsg4uDBYPgYbNwLQgQMP7M78Lfz75k+HZvPYxv
M9ivrm30GIJQDUiDUv5oT78aCpGDN6aqDZbDNhhTzSrj32tMon5UPI8I1w3c/Yy6
AB15UchjiW1gIDMfSXk1B5JNCi/gfIGhQH34V0QK6ibFrwJ+rl5gM4hCMpwR6hBh
ztKuhV5dgOkLE5ufamy5MpXX/i97UDQoJ+m3ApazLERHLHuXuEDzdWzSQbUCiME6
MJZuZbMmsP0wMkZdOln/t9KNNjcK/sCGaSvwNjewElX4qQPwWPWbCHGB3zCty0Rp
diNgfqSGErka++wrnGXomnVQBwjk9arJDOX6c1pwu0l+8lkjIovreJbBxPTAAPYf
5lZkQxgufikuLclA74y2i8TixKXX2Cbppp7qqLYTe8gcEgwEqIVYucV5t6f/lufc
5oLhgv5i0I5dYwmUavPyrTGeuYmW0s2QWN9xSAurR2XygUJV+TIvhVXgwTq999u1
6BuJqveTGKvtFXeajgPQhLU420c65o3utQikoJxUFcg7KWZWDXkdr0qKP0Zhib/p
n7NuB+iHjVxVco0RDtvHHP3grObbaJIlG5Ut/eee/LiikJomBedQYZbGLlILgj4k
qcXdDXte884NoTx3MpqJTE1brdtd2IjZQPF6B4fm4ZRtWpoXYYRxmypN2meZ8OO2
yWhjWWuRqsh+vkZAJlLHea6pQEbOU1J+Sv4NiPF2Cr62ADdLyv85JyNYUvpok8Ne
Eh4AY7B1185g417qj3Q5qPbhqUc+bk/slhh20cG/IkIJ+jwQzxYr4lvmUG3gHmb1
g531boICHEb0KujYLd02OtmhRxEuhIgGR1uT0depEOE7FAy4c2wmOPrb0qksa0eJ
KPIPh+RLB7SvSX2gcN7FON5foK55PtgNR+TS9eEoqNmVzVnV3WXpyjJ8FTq49x2y
AHEVdtluvOFtBeyGHcWa6+f8zJc2s13AggHIpBlTAer0gt/avCkffNJaNEnDXCPY
Kg0ZmopVOl8CF1lVMfYUEMIagULLOTIF5qv3Z7n/Br8012Z0tushy9ZTeUx/5NGC
OiPfPsMdU6dXECJ45Lu8PTBzga+W0SGyIoiLce6llJZXoncbe7P1ZNAfFKIyyjzy
alZrNfmO6JTXFMA5xsZ+1f89TYqN82A2mm613x5uY0yIJ7IEJGWSCRVIQAZ7Rmzr
YaLDk3BAkznH9X45F1/p+zJGTMdE2eD4VNZPz6b8Q4i3FssEK6Wg9LwxabyMDGiS
LkkIFsIgtAq3ybeNBSTrdMO55of7ZnbiZXsf2b/8zhcWALKBfpIyf5WbjX2A/IoD
c1QaMFU2PbXk6YJXsNbLEqNdd/fMaGbZxBiA40syR4zkLNifaAd1U6rgowe1zNRe
flYHusNAH60GvZxYL9EYD8Zh7dBNLvFLP2V/jwudgjBmuUrSw1ZyawogSEVwdMMW
/0z6JnuPbpb564iP8FZN20zQhI52sm7wVDd1pRta0wsBCJUdo2Z9em+i3boI+0dk
YdSJtmaQS9EssyeRiWXTJrTD3EQnwW+o2wsw3BZ7PhFJ/bVE6zvGwxMcsEeL/YCO
wz4Zl9zBp4B1V+IrHEqGHhJx8BbpV5m+T5dZ+lSl1QOa55weNdkom/onvBx3z3qD
Qap0I9/qJX/NeCJnm4opaC1925AHjDR1PaKNFRIDN0SQKFMgqOA0Jgvv/0ulU3uB
C8hOeDshiMK5qZ1Guz0EiKQ6kjS09fyHUiIsHx3wT2FELu8csjRn1PocX1wODQDF
5A9pUxXOt5h8FwyYLxqbzfzdhTD90B8zV55iYs6xPCfJRDjSxgqIPpudXIIdL8R7
gllDHptG2pQgFhwmc6gY51vUJjuxq6AkYtyXpMjyhRCzPbBlTsl/RS04BLKuqpaJ
1+az7FMksAezYIN4GqfCkbiQSUB4RAQFESblL5wKPo1040HsfEV0kGh6/mouovPL
3cDRfuK5hRnS//pdEDvQyCiEuIJ+PI+9IdPydSIpiqMzjaMshooUqEG2w2Ggm5It
jrcvmGUkbl5sh7dZ3lUA5dOFYtJ2zlrb4DgF6hxS6j0QU9NGPBcHI+ouZJuDqp3l
vYd4QsYO2yVek4M/PKsa+LUqvNg0W16Z+vYYGrJ80rNBDJGRhIc1MgUF9eXpNzYJ
+03R66NV4wx0IiRqzZKbXwsagszAbh01kc7XRiH5SPwJN4vSvdrtASy+j546zjd4
e6uHKLCzsPvACANlwRzpDX11rSA8kIxYhWppEJ933PUZFgV1NBkPENpBwiTAzU6L
OGRT9n05w0eoDdVOb0YS+q99inz9m3aIW0QFzVvv3MMDN5nzG0vDWhxUa4FiVsqB
sGm1pA1xZIJ8ExwJs6IGu8COxeIJnE3kSVFKF/G+eqZJJoyIskN7tOpOKAn6GLFP
3InzLzHoZC1mTknHVWtNohs+5dehMh8UGfma82XMoSaTV9IhIgOIrroP1rrf9qQ9
Z08H8GYIzwuMkYFmk+STrWTXl0fmV+wo8Ig0AHouBS2laRsdfnsLmxpZBcOIhdb1
otOgJsOoGkS/WRyVnrLTbUq+olCtDHfRZH5LE38C6rtIYQsPbiE+kxU1TdRQ0nV6
QFpmTGt11s2gGP4psAWyhfdFB3lROzneYyUYaRO2pCmBB9wYwZFbMOUBrl37H8/W
2sW9ZIXwiWkKaZ/JOfLoVgwa5IKkqJnhIuvujrYVeRuPGq0LpsIJU3OIag+LGOgz
Ljf0KuX1vBAOpkhQ+B1NwZQw3rExkqSOU2IL3XuvPecDeMALSor93S3i+yQ1SNXG
o+9ViD4Nj80lb4oTUPU+Ly/H7nq+Dud4TrFMHjn3Hj0J+4HxHWYxN5RvvhrW1eAW
ZM4SGmLeAEnYxaXPV3AdqGf6xdpKaCre7G78E8UfoH68k+fp/TRRIgBsS1b/B4P/
6UKp2Sge5FvLwxcgyGO4Rxq42y/Pp7CK56gLZz0ds7FbkT54rN5H0XcXukCohr3N
BDVK7EF8wxmATjXp3sCTcMQT0M7m1Ao7z+FKG9I6Az8AfwfS8uHMRcJYIPZo6jvk
P351ie/R8Rn4f7rMzg/TlUtkovxzmw4qY76tfzsvoaFLu6qpl2tb05nJMz/fll/Z
NodKeRfRPXNfich4NhuwJAAQ99Tg2PQT6ExrgfkuJQ7T/dlKjOu7MnTP4fNLu8qr
Xp5wZZZ1BN7Ew7xyxU7vcdv5uGJa2vmzri0NPhibeNttAg+bw12C5t78X83FMatz
rgNPlG1gdITH9Y+1K/ZtG+q49IWb5NyLZr2g00cgmILaVzEf7yAuBsJvrRXCPm09
rEEXspHI5+OFkdHdIXofpNRm7L/Pb9GfBvCjecuZSYfGI4yF/HUdhn3RxTzILjxw
fQZCQ+UdWA9om2hDpphRi5PCzGZFzncnEcU3jr1IltJmlPT2wbVuUu96tITgfyxr
m60JYrZl3BafJRuE1jAw2kF4PSb16wweLAWDYKzw0KYtS/UM+9Zo/hwyUFnrEQvV
/s7IkX71KGIaXXizhITKXlk2ik51FuxIPFGisqPW+Y2mWR8M09h1IdNlsa8Zh+0K
9mn46Td6eX0b0xpYztPChI3lOwilsHUkCLYQoM+YwQ+F6OST0VXSqngnrorrGyCE
2bMWB7Njb3ziLXznruvBpVfMsOCqaXIDBdcJa1D5fsqKSVZEz9/TlkkzHnb173Wl
6EawzaMUhkO9XqPl2H0sldBt6SdVwcLIf0tZfsRtr6s+BRdcCYiY7g9BdzhewfRV
YkbDdkwL0/InicoQje2GCMXnw/o7s/926MSEjJTRx4mM91UtCJfCkjQ9x3jVKE/w
9T7uouGg8thPUiXEaHUF8epr4SiP98Ji4w5ZI9oUZ1W9ZT+RfYE5rXUjIsJpbtRM
sEuOyd5TRMCESqT4k55+6s6xQcyYtEO15cqJqHJrNKomgK19F86rVDQeRj7ZtLWz
WHmsKTmvNsMznaSKY1Lombsq/xA+U7afMXXO6/9ytk8LCIAGO5ZWB8POyltvoyau
Y66cXjypSB3CbRzdMFGQ+BeWCWsRpFovr01VWkNiA23/HQrIpg+qPEOKKov38GfT
zhTtEY4rRc3e/4NtN9w8QRrUtugPpLgtiBeYt9yyGE7u5CHic8JupxRI2LoMUdU+
NkK8WCPsmn/8KYbdjlDsQd9QYHJNcWyjsLVKpZTPjeswuXnFvi6Mb4Oq+2ID+iPF
pxgFL6yQrU3V+7nwKN/K4+bFsp/pnijoGCcRt7nYsZIK/ULTkTbyjD6ul4yUyVNz
xcjrfNgU8KniNlubfzxhJnLpesew3OBOF5V2UujE+WpIn/gLDzsguXXAULfhgfTH
rKlLx3XxyexH3eJJZcI64D4o/2O2wbxSyIm9yfRctHTiVtXGE/sSZerhCF0kHtWi
EEcj0m1OsbBKNwfTjmaYzLgc9QRUkbNbZZGN4jkY4QhcXMEvshaP3KDsRl743dk9
pnmYHGuj6IcUJHKDrP8W12nC9/AIM13CqGymEa1KxIiOyLRG7kMVMEhi/bnCMv4F
cPdHjHPkFz8w2fW/cqeJhOsgA1vOp3Pfetcs4gpvReWRuMw4VIQx7Q87pzDuvthN
Dy4jtxkY6vQxDqu33msfne8vP3AUU/5nKuO/n1xXZCoTbRuF+v0qRybSHmgf0KEH
NDdpyfUDjr9hwbQyLuAn0svWd5j4kefM0f337JN2RquaxxrLKdpBSc4BNaEw1WKg
NiZYB5i7zpv3JLx9NuR2XzGZpmcT/152xiAfmGvtJ+EXifDkLnFjzZZuc9Solak0
8Nkm5HtWRSgRhfDW2nYOKtsJoTxB1maZa+21ADrRVRXFt/B249H4UhnoQ4ZotvHx
uRPNFPAxGdfvBa+gBpvi8yTcdvdAocL2b+u9jiGbdX9ekAmCjkKM7mFik1JJaRmx
+vY9BxX/xm2gxMMahL7jxzWTIyicKMVJCOZflkreKXrT9lAOoVJx/APsYEw8aEF0
22vGKGyIiMiDmLaczpC+E+egFoVBScAdmkYsqTa7vHxhbt1XKWmS2s0aFZbLFfCZ
52kpIbxLbJpWONTEc4u0eJ8oIbYP/MWS3RsWcpBDzZfgTsAkrPfqGauDI5dehTN7
jVCKBTry9/93a58bTf9ZaONHzh141TW1qiQ0wz/016iud0pKzsr/wm4BFgjoQBYy
XLgA8hgl+0ClFKSs4NTB2yXjuWWHg0h5IryBfeXNq20GlHBXJv3AG7blHkCCT3v9
paXkXUZOb3WxPWLVJYl+KwbgzxgZkqxFmtG3nK8QVOwm9vYpBkQryRi621cMjFa/
e/4WLX286HT6PXuQj4OehnF8wAjSUy9ASkSmJoQ4EmUak+kBjidLWgHTd9DRGZ9w
grSCPKeH26MwH1RNVUwvd+eb4NaMIb6+op5br4G2/Fw96JrPmpokfGyaEf9WVgKG
lOzkQu/5A9ZN+tpoHVBM+yw6q4M3SAeLrpA8baN87hG4lHT5qxW3o/dUZn8XrlPQ
rQkcfyfF3NiP0CHj/8jVa34PLTnSecOmVR2B0puwFX0avJAR07m5Jk3lmIdyxR0q
u5S8k21CY1r/uF2yh6Mzw1Mw3vW/qvUoWEUn7CMelNeGlePNnnqXmB4UDDSdMsBN
hYH6GJjavBxRg6XSyY7HRKas+J0M4yZxF9xt/MvzBmuv/0FS+gV9zIl1Nmu1T9Sb
Vbg2GRnq1HvFgzN9QmwWvJRgLL8guIMNuoxDU+inal3o7UJIrGbIo8XSkfGneWqA
DrSwDyITXuyMq96tYOodSw9ATHQi3ZvaDFHqtht4QadPdXA6GFELDJ6AfsgxZ2ry
AaoQoFz8j7JIlNVObN/k8uN6POXpAm+0bJ6VuwimlKMmiQVUF5gyb3BwdexZwCVK
Nk7zG5pm0WrpNfZfu6dhuSFjrpb/Kvqme9DH+BkYZlSQJdJbeqpb6sATG+FKB2fV
1AgdiRurOq2bAX85dj/LaBHO7I81RrNQw05OO6VPCNYzugSV15SSxCy8ZdGuk6/m
30/jsxjCa/kS6XH6mOP4RevVbBeytC9UAh43j552l7ZnW9rghSJfShMNEQOer3pf
UWWhnUUPZb4f7BShISCn3QWKePwp59kibV5PVCf2wwId51ByUImTQx3K6Qq5VVLT
dlONaLP1oMi6rIfWpekHgEAJJIaxPZGNlh5Bq9qfZ1Wt8NbVu99LMMLnj5ijdzMd
9vzOHpExnaPDXOS0c5RMxMYfAfF0W/rN2N54GJ1KXEUaAc0GwYIGg/Uar8rfdW6i
zQD/UdIefRF83UEmap+rcw4H3GYdD111qvPwjeWz/jAEfAxixGf2sT8J0hE09x+q
aqgBJOqZdad1ShyWvQYbBd2pLcs8anu6SlrLjAP+VmlRZNHTZplxGOCfXB0p0u4s
uDa77IIoPDRJ5PLwSv4NkFVAWqzb4RfhhNcWLzDvjZh7q8c0py+yx8z82jnBwyjg
zCjdlLfQW+KJQ5HrAb2+FuNacajjuk1LM8EWMV32isdXCafYSBfoSfOZ+pckNTMl
owjm6qXOXpppRuDgMg9GoTvhlljWXe5UayL3HBoiJAx+9flLg34bJ1aYtlZ2ouCa
1Nenq7oNEJxlXNjHlUFMUEa/eyR1Pctfjx26TODzJ94cDDo0uRlNsH5aLnDWFudF
qOG+UxAUocmW6g7v7Wr3uO8hQV09g2zIHTEAJlVJef/CeUzfWXkxobnHHvnACgmf
KHAAp2/XS7teACTJXoNQajmDLuR1SkI+G+Ysu68T4BqJqZIkm8LlvlUQFJ0AVziP
dTnzYjqdzDs4wsiWOdw039/2UU2/uiuSS53cVDrMUR8fzLtVqU8qVuzE8KzzlxrF
xNvFy7Sco7arjluXzUsv+CjfddsD3gq7A2poelFousb/I3WpWO8xJHRP6d7aSUFa
a9WFACViM/T9lnzUL0Ifvt1ZCXEOeJA1GZ13bRUZdA8WYBhDlt/WyEtg0hLI54BT
5GAR/bt70DR/Cl/29hjYJOrK4RIKXAICKjEVXm/dqHM88M+ToVH0G1PWd4XRIwFf
tLrQ2foKYiESGU61o5QFi3Cr8FCACAqi5zwkBt3tFYhpmrPH+L58ZRR+BpiiDYZa
huhW/bNMHJrAdKBkIL/HdiMDNw6R6gCdQ6qXURB/iqpnB4RpVBr9/ZB/tzIqkwEE
52DxGYJReT2x0tyfvdJBhlm39ufpq+R6YNPQHmS7D/MQKbLI4P3eQGfA4HheggYP
+LbEHT3jb7oFCmcLlyGxKqe9AgZnu/9IUCM5JMiSBmlp87EhLXfJIUSCTyTO8xuw
rg7uV24I+0RaC+CMKIxJ4zr6Jh/D5PbeX/SFDzHA1/sCBX0tz0923N2+GvWmWzSD
5YJqXu6kElLuJKP+pJntlIM0e5xA4eOC8HNzTHYMIoLMXouiS1RWHWsK64DUhSfG
nHp7368lsUpIPZPwGZuzbsBpn9GMr1BIesDpTMAwtw91a/lmCPUktPXIPB+lAJ+6
Tz0a58SSgvO4ywW0uMszVI7k3YtglV94y6z2fzLApeSgyC1r3T9LDIoss0JXKbuz
gf7QIB/U9uZOvtuFz2dRKFnOqhEQj3ABGweP1WCzE8keXIBrAowNTYeMk0V4qQ0q
PJvFY4lsZIltN2AWGZi2dcXZ4t9Yvgj+FxwB273upOYFylVQpB62/bK5Ga6VrEYC
fA+IKazflcibtGTUEe+VXDRXpMffGz02nNfy//NNHy9NZl/4ctkvj/4hrJAjgiBt
zTaANVYnGxpSLS0mqRZB4bI9bVAYpl8cGt1551RFGVMUGmD6I752cWTajMPs7gPo
c/vJ1ZcyrBnI6CtJ0/IBURHeaYyf+OL+wvj2lWTOsHUpCV/bXtNwyih4dSB6viKd
8F7gli7TwBmO2pNZQ1g9yNlBRRoZ8MHEw4tg6bka1qG+UiQE1EQBu2OxVjQnPHLj
JjNxUTPC4Iem+OKlKTupOcmzXGSmUVVUiVmC6nQpbh3KF15uDTPH7vgHbb1NjwGo
kuHKokzqLFrvh4Y94L263YEopEDxDwU7lGco6Ewsdmc9Ma8xG8FtR7Qu2ZgpB48W
hr24YX4dF6FgSRcBnBh5MYek47kVEgXzPazYu1lWiDw057xm64f1/NvMQYWvjUdQ
q8TJ6IBE7z6XxO65FAkDVUkrpUQbRV+ngjB0wxWHje6aPHgUdNVHCFOXiJf2yVbu
ASOJ/Pix589F273M1pheE7zptKe7Ed2rLtnZdxNoIx9yHkzs19/gHXXaCobuQcjU
r+JFcRR6MvJinrJI7G1gsLVBkJFpddGNh3OQcFYBquaEOaQ9XnBDDYruWJgeIlvi
Kk/X5y4h10JhzyyAQvJyYK7Uf2ayaHRRjfEB+4prDH68jU7V1gdfiu5ip3KSQHNH
dURShMXG0oaKhMPkaFt82bNIhE2VWJAzjW2M997Rk8OHAzul3E1X1yqeoKfEJUUD
HVnNEXloJ9BzyEFr2oksVQ7jFehlLTJ7nytyNzJ4WQKxBlOcVay3Rt/HA4wCrKXg
5JfVC2OIQPb3kbZokQ7ifmJUO1oLtpcnHYdOn1z3uJDARp9oVVNumkrza9LvWF3b
NJgjYT6YXTW9S2iyX4oJy6Y8buX5nB+fgj4KhoK6nDpkfUnBr+YNQ+4EvhKvW8h6
GfK5+XDiIiQEYWTNTZK2U1mPhKTzjH0+BRAEeuOjcmrc9o6zdOpaGRKIsWutiICl
zm9ccxVaEX18KXjwoQ1RC1YVRngDk0HniuSrrMjtg624bxihbmDcQ0mft1nFJh0f
sQ0l1nr9m1NuaNXnFx/nAommanJDGGw9hFXfzSjHU7XtUZaD8FvJdoF1Xdg2/5dp
Qa1rS89p4AMcrGjc1Xxk54KTE8pUfFjPXRg2p40lRVmgIGF1mJ1R+M8zWbtA6Xgb
G3YL84HK01Wqyv8NiBLtUTfLJ9yBngbnfCjZ7Ud7AJbIglZHKX2kcSh6j0lqZ21d
3+t7rBEgIEWw6dInwZYDD4RJ7lJslX2qpSziLTLn89pIwqHBfeVdMUuv61wLZMDM
oMdI5+jC7MqSI9fJ5wV7aUtWI2IMYlZMMnffYuhUZClWYT1t7uUcjZqJE8sinp33
LTzttTBvADTV5Rd5Gf1XXuPsjpKSJqmA0uiAOGgFY+cP4/v07/I23BtQ6aoB051H
cOg6yatlMnpTrbgc2gm3UWcPxvSZEaOO0FRnl1PIRZSNZQEUEKN4XpR3J08yO5bX
+6Of77l/0DO4BtOD8DQyCqyuHQq0fUVo42TeXxCSVuZf5/I1Ca83HK8nV3NC60fy
6kQAA0vP+Fn2vj3bxv6JGxGFRymB6nUoPZbjy6f2WtWV+vuwLGXntYuznRYMk1KO
dI0iLZXkqtNdeB3M02kVfV/YaK+qmaXgMjC2I1REzFthAFM5f9BS83o9hBIrgxXz
8tmBwVGtBzVT1Qn8qOjn3xCxu2Rp6A4HF5Z7tpnaBOYm8ghwBQgDrfwFcSLojE5X
KWS5HihCxJDNYv/XA3ZsLepC1Bj0Ux8VJeY/z1/0SOW8EWBXYbQL3sANntecLFMN
ialXlnpT7Dfu9Rl0lXgUPASUxSEIhwshaQolj4SRSUp1c+4/r/Oe4O4pm3yuo42n
yhZKPK5+NiAac7HDNhj6m0TU9yK8+hK9WesWs1Ybr+ihVyYakZjN8g9ZbzNrhxgh
f/Vp8a7KFkZTsmlc+CJpozqoNzLF9NXs4oB2Cx4C3802AJNq3bQRy+mwv/m5vzri
dRj3MrvzSzc4tSV/R286xYz3l2gkhjIOsLpMOZv1wVsc7sq+rnnFnojZWYEUAUK7
XUIJd9CvNg9CU4Pzd4kNDYAx3zB4PtbnXsSlKvd2r8iTScvJA6CcPHalp+TyFbEJ
Vs12D4iLAN+Dscgj1CvyN4LNjLOEP4uZ43q/AXmKuKrusZpmpE7U88I6GGl6Ezn2
UI3QOfT7VkqF0sKOQaqRG4NBeJx63cT2py4yX2SKaoDNJ6Wf8B9QJXNoXlPzlN+p
bY+ML8a5T4kVRoVYRn652Ky7sowMIU/DmZ23Q8NscqaF+P2UE/G9FvwH5/KYqmhA
y8mcVQe3PsawUY56ldoAR024MeF1nld0sjWYQSaR/kQLsL5q3YW+EHeYmvoYKTW/
vlEXxkHK8Qo8PZnup5o/6ojJs4x7qa85zRk4Xgz4CIto9+gQ/HMTwIz3h4Kt+Cu5
ie2KZRXOZ/VDA/3apXZkln3mETHw1SQcMj52PnU77bH76vPcyE8vHsoHK+WX7yg5
72XMQm3xjDEtwCN9MrT5c782UKRIbK89yGskx6b2k1aVblTHi24UIFBNUJQjmf+3
zX1bpy1EQuCx2smD7FSN8tNyQKpgWqpELiAXGNz1UrA26834xBF08v18ifJv+KRE
B4EXB0AwLY/DTiFRVJNS5YAoZtynS0LZMHDn89p+BMX6C2kmXCTDrFUy7+wSH7Xq
HKFkX2oxClkEZV+CmICaDb5ZcgOvggXhiuKqC41UWKvFTi7p+wngtS98Wr6DM5Ev
hH1/1Y/lafCaCj40uuVohx7oPGcOj8mcS4aHw62i7UI1CWBl3BfWZBIXudJwew2m
GNkGZRXs+1oiGiEgZVgnUpYtIvYUxDBCydJ3hhWHBNOVURYUa9cQX+VNe0KPzO0z
ov8RqOehdz6zCWwmLmz3n065NLOdpXBDGmgmHFEOAQjg3UfebGKorq6wKXyBMHDp
CxZ4XMNWD+r6BAqos0k2rwPE3ygkiMMum/lGkUZopke+ENPHq7y8B9dZwQlHaE3e
OLp3WP32SqK7Sq3AhFeW6Y5axf/pFiqECdE6ZlJUmO/hxCTPr/VakKcJl3uozn7L
Pf71+5kjl46QZAVIP46mJgfWOaOTD/QW23t2co6ja4joLzyGDfq2yleRqVjzE/sd
DhA86W/L7/KzFEOIWRDALAs2GSJRZTuVCf26J2P6ilgmLF/sSy0mng9js0QB4Eim
Hh8sOSb8w9rwPUYU1nQM3oPGkbSVCm8sVfYpF7IATRPdeuMfh6HIrkMS7IxaFEKd
QEg7WKYAHYs5Jroisxy43EczP8Xk4nSGbyyo7xa77zgJzQABrcMa1iBTfoetONkP
P46vhBOnsZtiWh1omZQ4GWwLmrjKoTFoHu210VxEQdnisNiyzDAInod7jHnCFu1k
dgYlYsEoLWU+ECBuPfjSjzKTUfZUsmACaBqbRycRb+xS7Eg1fSthTMDiRka/Tk7i
59fLnmiZFs34T/Wb6PPoB79bF+oC9g8VsxZWvh3QoIwxqRynq6OELS6d84jRU0Sn
yooho9AXZKqF4qTzNfyxdCWqcGzau3gHMlpl8y/KJ+eckZ+Q0XMZK0vJho5JAAgX
zcVUI/bhU3+Kxp0vwntBT1F2obEYfiBwDYCBzpKBbsV4ge8rnSl4gYecyHJCKr/K
aQio3DazRneZwR7RjMjJG0RC1SIwoYrVnNO2SDH3u0kpAseT6Tq1dMBTtguEvLzS
uiouk4CasN6jhEEg9UU0vGFXZDlwSDgTCUxNrHIiJq+51q/7Q3oBOnNlV3XPkMaO
Tmj0XKpA9C4YNHDWxJTpx+qNc0Lz6WZSTYCUwKKwbhrN9UPSzYAyHC5xB0cDkwwQ
w/XyUq5EpeDpwKEZaDfsiau+eP/KKHGqElsPqRMdb+3ZZmMzAAih2fsHv65sJAuq
lsyBX9hhM/aLK9zrqR2EqSwEhfhP/riAX/VD0+ZWd4eiUW7nPvuE5HZ8SMKTpj/b
CK6ZnD8whiuHkXAE/8a1nDUs3KBiYcqg19oVQub15hGC/ynJ8iChpUFMJp3nyecH
coqB1WJSMbxufU7GIqjERV7EbZ2BTgH22DX8O7bfp5NafMpI8/njKdqvsqnScls7
bY0w5MNQpgrUCN2NUtQSPgOcJwONjC1B9egRhfNDefjvLgqfj6WW0nRPuMrb7o+L
IlFhya8y926DhlHycbKw/OWyXGGvZfY09y5W2ygu1Bn7jFobEtY2BlCj6xGkdqO8
nZjifl7WZfuYzzd7ePgc3vpkAF6e1JRRtXAFSdcvsWlmtcoKQuHbo5Hf+AuFR1Ek
DzRahqzHWGn15HYoxI5pL/PykM0eY9JvmC07ORrhXQy2VGYz1dq/PMw4ND/zOivc
4hgey/aPgtC+7iK5OYW9n81SKxwQ9VSFRShjImJQjuiT7nQG/loeCxGYcWyW2/C/
MW+Px5ORTg5X1kVhEBbKLecszpqwp29TOjBm5R7GR9G/G4kdy5jRl9JDSqR0wkc0
d2Vg7k/7tEIKqFkColGtBYDxJQBlaOMarvycbWuvGkg3boQT2VWNunNpe94vI+Aj
V8db2gEN1me+k6vRjZJEBlqLQYAZReO7zVwHTgwYvMPYwcWEXTwigbL/zCxGCNiP
3BBI+/BNtbaJ3mmj3NzadxO9qhkNdonpijTsCNPFdymESVcylUk671GmvWwK3iXc
D4ulaTq3QzSHQy+l3jmBOUIQizQZb3R+f7rPge+jgFz8VjRjoU7EVhXso1xqp93b
hVBd7L+0NyQm2PtDX2MS61MNLekkx+dK3XM3SLB58xA/7XWWoic7x2kHhqxx+6k+
S4KnsX83EwRa5FwNeOa8FF9cgpiBuWs2JUvcP495ZWljIvZB40uSVDvWVpNeg6Op
GxyCXoJV0jD7dJyvrNxYAh0fr4VfGOiFGv3RgQ3JlbeE9RKUvl+UsFmYpwF3bGAl
DLxROHxjAmWqUD3lLEFl5iQ02ZF2MRC3Uvt/fDyem5dOGAkMufNUo3MMT223GwQj
YbYADYjmbbOFpcizzg6G0D/bm0tUcRjXb8HjbFmIUZ3GZZduj81IJSdZROPn9+3I
zS4kOC43srFv4SeuisSOSNOI8uU7BLT8FvCkYSKNYvHdVowGnntG7pmawR8jFmbe
BdnxNsTNSKkPX53NBGBzbyldNKiAovg7Y07E546gpFEWXMWoCuH2mBFcAzyRGqi3
f7E1n8zxsrw1YWP35CqzZoTXJLsH1Tl3MV09EJVb/NMrrx/woaG72jYEADMJkgg4
2JqBw62bFiR/7VC0gArxE/ff0Qa45EmIgi8JzELG9QuTNagZemtwLZwtGNBHmDKU
crFNGJuo1pbwBvjooiJ9EhsGxjO7zh2P4GStnBiHk53xzxv3iJ1BL6pevhPJOfRx
Zs0YEfv550sgORyUQXyBt5CnjkD+Ean+GZ10IIfxk3zcudpHW6QLO08oUmsObtLW
Ua7on7dHlkxKFsbduMn+qgkoF+KhBxZ6k3rcpl/hqtBQqJ6M4dhVOBpkKbGQbpCj
ZhUda3Hk+IcEg9thbcJuIpZ4vzeR7sLFnk2z5OJFsfL6IcMfTNGYO0MjPGvQMQp+
wA6htv4eAxWMbnx/7UjvvmZQUAQuGgFW72Gd3cGMeglMZUfjjjjm2VViOnbKe/ab
RGqnfN6gThoZ8krDmQhhy8TJJv8q9+x6XhUFyKJShUvRRpndSSSUHTaAY7oGIiPN
wODHEl78uWWEIsihknqbw186DU//BRg/EOX2xQchmSvwUkvBwPr/NMTRQXM+h0Zx
NWFhxH7gchuBaa3dqN5S7oZizKrxnxqomuCdmIEDULEo3KA6Q5TIo1eIpyq+1n8g
FRoXsIsCnvI0U8U946D1rLXS+UdoI0JEjPmFHkGEoVl10+UP/3TKsAkzc/zsGtzU
I9HIHliEboPlUg9CEDFFKiNpzfhtF0mexa2vOcH+jCihDuGlG4D3/U2rqzVfCvOh
hBpOqQswQcAVpd0Ahi6aaROEUq9skIRry0ahujnTtEBNoTaPVyWl1Clw5PUA/esv
cWXK03NQCoMgjsaruIzpNKgUZ8diLIF22juoFLUK9JfWjP5MWFWZqnYdWCAOEc+n
bWtHYA2K3GDdgGco6to5/pTtHiMVv89BtIrVgZ9AFco7m3ffVH74so2CcL86D7Cu
qnrbHms7ijGJZi4XT6GMLiWs6mk9+sL6Ez+bHM4hqqe5gX8HckvEeKnSE31it1ui
B8IVwAaIGBeMhpZaJ8zLCnjTbM0bF9jWcfWEOvdmdC+18bU58Rq8lwFLoasweQB2
FtNhkEbSwxdWhRxoFe7hiyoaY5AwN313MYuYoUF74K+CcpwKEglYOL6R0pkUwhCn
k/CQT0ZCFjuL9C9OpDYkESl3DsUlQ5I03yvHFVaJoFB9IBhsDp0F6YdTACWNa/Jw
3B7NIejDNArLUEqwdfV/rw1LBSM/YEvJdll1i1uGRqQ9ulxcS0V2OHJ+8dV55Sem
4c0L6/kD5YPiZVxfjXbTxiBkSKH3eDNoZfOfFc0MiHHLh51wbMtLCFY0cxSFiVJw
rt3E9LUq7vUG4modzLpGqhnK22jdQV1cb/EYgnV4wlZ1IXMLB/sz0rLXZ27SCt0T
PcLkP83Ptpo+Xs/lGE7Fb1nVSK4AsJnIPFjkJJxr9KDw3BLbLqktKRxR4baIEGrj
ylprJ5l9/yoH6RMC5qG1nKJJC5CfqdWxZRN0YC9PwE+tS1Gd9dPd0sm6by7jj0yi
pPypJaeaeC6IeJjKAewc+gyCUuhM3Y9Z4E/32+VfdxT109YGAW7FhbmEU95Lr2La
gIfMGzIBTYDO8SUVfePQ4R8XQjadPraGDkTRgtks+fDF4JyxdAABH3jjf6c2u1DG
/HmEdQJdKq+cT/7d0im/1/T5XuEdtVH5ahaeACeNOKmvNj7r8tRalvt1MbgdxIK/
IzQ5PVOtb/yyTuAhiU87lH5jM63C9XTfauh/Badvyv0m0ga2/VVzPQFm9u5Rlqr5
K1ENvuBK/rOCk2dhKf+Cp/6w6RVOeZDAEkG7JNiexKZ8G4TWDtUtwixiMESjP2eH
C3ibRysMjTfzBYMUljroX18RkxyWybIrVmToXOzLwAosUsESDZ+QnKL+wM18+6Z9
rn6OdkJYdC4D3A9HGNwmzNlwMPfZZM/8NxRdCHzTjxVN2aJ6F0R4mH3uBqdrLfLz
ABE/0xTv6y9ZIszv29ganLaYGvtUy+s86N5SD/hVXHBMl1moUQjuX98YLLFhUBT/
rmRwGlQ8tbldImGNDgWGCe/06Zg7HEEymiICMLXFLM3lQJaITkHkK3qFIbTXHXIq
OmFMouU5k1DQt7PhaYF+AZpT0o+3kE76iJNLu+iQtRHsLdkkMlxuqxt6B8SFJXTu
OZ7spjzA7uK7VPh5uOrJjU0X7os4dic1ydK/h88j196Ng9/oVBlBtLUzwpFSTEuL
Ft1QaWleoIJc5Di8b2bp5C/1ydDQmAaws/b4dsLiteuiMbE+RxoPHMapuLL6CF0+
kNbTMhb7K17nKlea2U6YwcV72eMF0SQUxVc5xCxJ7NFgEg6MOZijhgv8O7r3D+nM
hi/DXRyGjXnl3LxMyUy2jHXMS5hX3FZsN0a8A9E6B+faSnOYVurp4giqkIf5QyaI
IpNp8uNsytahraic3iwUt2a5GQXh8CkINPozpYleCE+7IVadtmKmKKJLAFDPEJd+
hyrhubsbycCzorO6QvzQwmNzj0gCPOpYPh5ySxcDzz3eUqeV2pZeIIpGs7/pnRq7
KsaBxRV4DGIUaVwVCQF6ZFf+hcgv0yUX0kuv8KgTZ9LxuSeXYEm64vtVjW/WYBk2
p9W9YXvmG29rJvqIv1Rk9sHP2IfJgposD1RVj81Ps63oJzlSq5lxdKWu3h9K/sV6
n2byp79hkr2xoL7FKl2vedzW9XyXw4x+rMV/9I9kXS2sd5niOHRuTAbnAxD3/RlA
KRRUnviZWBl1y1Fn+EAxDM4tDyGsl3g+tE6I7TtqJ/gk1reCm5o8QSsnCAWLEqAl
y2UmseJ5yXGTplNhABVXIZ4CmsNHkTsJfzJi089BqKuuLbAMoTwRCZG0MR37yqia
6iMJQnte+KDMHs5qu20XLnDKu1cqUQXUy3Cmso/1NVjWQ12fSzkadAAIIgmuGVJo
W6dqyM7x7WAn6sqqCZGzefZNe0Gm9Vj8rUWxcEXMeogtjPxxm25ju6wlGfudA8Nj
nxgk4bbaKbekJa+uDlyRIwdouHrk/C4Itafrnfaapv94lRxNyo41c4pMtiYEDCzo
INFFkprXKnX0WuLFa5RhHdI2EJMvygRePxWuuThQKJUCJSHCukPRAv/bwNwuMziU
KR3rjJtaqdYQhNJz8w8QrVCAiiWL+qi5bHAdR/JzxPqem/QuNXz+L/7baGV3mBBI
28LIG9rUPSMjJXJpPHBSZ+oc1KgQP/ghS1qkr8MBOee0EuOEHU2q3Qx1eqdvkJlH
yadaZAul+X4wefRcbtBye/jwngIxBv+hhheztYSq5EsHDjUL2nenSp09dBjLWznM
0GWmeaGRR32F5MldwicMXNYV7bD07bwfAPYvsO6niBVYV40ebqV3WbeLIsXGI3QJ
BTe8He92JiXvQIkjy9w7P5u57yNqfUVLAqETGzNxUAghg0WZK8rvSSId3Uc5YgCK
evJZXpowU4OTP3DFeuf2awtdhxPDbEFe+i1E8LOryPv6hO+JKmP5twJU7CnMY8x9
sel7mO4nHtbeeYt7QU5/ml3/nmgAUYQubEHxdNe5aS5QgUu3Pa+A68EDkmZ6oYBb
uq460Gj/MRP7TdlknC79mDTXPELZDdcQoMCGlM4gEZRXoXx1CPtDBUw7jF7SeZtS
JS1Mqxg4Q5GdL6k/UfHPNy3HJ4qX2Vf9axXun4M8TQOHPFKrydtdfqfswUkUlT/c
KLRrnZH33TtSIhB+nFkM95BoPozyKwTN7Rl+6YeMJsX9T4mEGx0DVUA3vULhd8qh
gJwibe570zT/EJtAk9Z11oBXOd42LIjrmZM7ALjYhPCbAIZ/JcJqMk9SkS/gAcUY
ofjU2Olx7nJCs9jxBkYFjE1IpGl+8xADmB8MpwHi8+tlczYP+poBl+aEpEfCIF5L
ib5uGjbod8L2Yz6b5nEbaMcehe7OAgH4pxJw3PxjBEd8OSBis9718RjSDijopNAU
C6wc8yWc86gMloyGWVc68uqWrEoeXH78H90zYmH7w2RNTvn3nnBYDGNGSAL9gAgp
tzzKLZkS/5K9MZTwFqEtCOM6fiMLOy/gvVoFfUi+KUk2apPZqExEvGGuz93kQW+j
8dblEBy4nB3/URVSxxM6BdQ1baQcfaXgwrH8iAZgf3NA1oCCQRZdEFES1GBdvDsv
On/dv514Lsmy41T7xWA9nmNVakPa8T1SYksjWfDj57QGHHjcn/6VuCMbL2wWQtaY
h1Gp7u1klR0cXPY+e9AicVbe7rmN0aP872XiuvjA2oT1U1/0MzvJcYeodAQjLhcq
DG0iCIc12uJXYmiAK7EnxkzQ0jrR+r3O8NWquAYVdxL2J6El+dyQvcTVlXtRobDI
G5TWz+KCiZ+WLGjma64I+pRG5Ujh+yLuftbOhg2wYYYP3v7Qk+TE6bXH9A/ffpF6
T5++7jy9w1U7J56a9NJtA4+NAIn694ekAoq4HD1p6y6wM8eJImbso6pvMWem0nee
EnZ/GfZST4YhYAn2KuhP6LPGukScV9Qhh73/6EyulARXg4q84Fjiw+BTkwLOdXi3
8ZscarlaFNRkGM0JnyCspYpJOD+7LLXGmZX4GlzuZuzfnwench3isuZLFywuyCyQ
t0brp2JH1jamVbn3OWAR+kLsBzwBQXpeu7rvZLCaMEQW/ppH1JVBOFhieYTqvGLk
M4o1ca7P3bHdFDOd+z6l0metKqxPuj63XzKh7f5u929yOxERnpSEpiVB6/YPkj1m
`pragma protect end_protected

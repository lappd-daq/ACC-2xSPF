// Copyright (C) 2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std
// ALTERA_TIMESTAMP:Thu Sep 13 06:32:39 PDT 2018
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
SI591/fNrjnZ7bl+923bKTPUVvWYDyrWBhuGI+pqd40iTGiAjjMh46uGa54dU07y
gzZ7BIM3Bnjo8K9/vjw7vrBIjsLX+NOpBojRcbs69TKinAEkaUZL6pH1cZNvPOqw
JrL1LtJ1mIC4k99R73HZBTPLPppu3eQ7xK3xWu/8+RQ=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 57744)
5zxcN+3qJg+udlAzqtVBqyC5aIFEbD5kDApn6ifXOMMdUyHEH2FFr9GHuKwwkKA4
llCD8/21MDYPx8mlv+9661U1cKMYCFzfsc+GhGLPFqQTSqk9E1isZqjLGx/dJyRG
hDrBEz2AQSDAiBO8BuBj4xzR68sP3xbPnYZckSJU3NRUnfK2vxzjALAmohUf1Us6
JTUWTirdNl1q0gvMdW4G7K0g0xrT/cQp2kjZfqHGkuVAcrtR+K4+FALVS3c2QTF3
uIj9P+emGUFi4JVjuWttPo8Hz8PQTwQrN5qpfdig6VpBk91z5yy+cx5vvN57oxG4
fQiQK+/xhXoNb/7ZNaYFqa11A5kiBgeS+7dyH9FmzPnDEPSv+3s8QR7bAqtG3PKT
MrDgn4iLYUy0h0BhDII0iLbsWNyeklPFXvDxAV2sBWmIcfhDLRsiopEptbpBXXlN
rHHToCru2Ed7wN7H4O4GS0fB4sK75IjphCZP6Z87JQupzzONl3MPejBSx8P2Z8y2
vUzz7kD+TwfbXBllL8wQKhtyXnCwOWVtp4hI2XiodJopeySRotNV3wlaq8KF6QsZ
MjFmAzDKgdfhKx2t9hJ9Qpr3jIjvBeelmiFbcvg1ydrAu27LpDHyQr86gfmGgqfk
SDDPhqorjYzdioeHeFEXV1HDyiaNDHpmhfV41rqu/f/ailkHfu8uPrP+VG51GMYZ
q8Q2noOpTjxHsCkU+R64CG+GMBQWNN4sSm2D6eDhZiLMci2KuQ0hj+chvl7nEzek
NsVach0dwF4gsUXa3ftPTMuJnZu1OxAxYuktogNwu2yeoomDBCw/C6e/ZkPorvva
bXpUJA8ARJ52Mt8KCtJqsAu+9xL/oyLRnPKsk43vyr8wFCDY/fmVT1pOyWk8Jmcr
Jva3KG8RWjS3tIxAMdrEYcDLg4PcBkDyaecD2irCCgJ27x6yxrnI9jJgSKIhU5z0
zFNrDf+DWqVJZExSuvET3gkEA6KgE4G1jXGTqyx7cxW2DLoJZsKb+LF6ZmhznFWd
MR0A0f5BGFYOdh+QXZCy+EcnPzpKR8cM1Txmh3jqkWaWFXw7T+rjDgYWFFKkf6pw
JVIufrSSFliYgdPGBmrr7R0OvPcUj/ZHAqSysHOwLBmhxXJ3Ozu8hy49tDT2EL3V
47rw0d2WkDB0hzU+BYHvSt5P/f+ctjtE8wEJ2sc9J26EZXJAYnLd/ng8Iv7Q2Dit
ASPN77xPi+WYPhz19g8uy6ltIOLLOyBpC1cLqkKT48Is8sByoWOfalHEiPowoMkt
BE4DLvGwzt8yiVLyRKN9JMU7ekRTmrQ+97okiw+Le3WG7tcDN6u02keGbNf+Y6eO
8kkEA3VY5/UgfXoAhW8/pffXizLCUpEYZJ5Ip4bMnrogz7I2LNHGujHmUb9og/7U
bjzSO5xBAg/R00nTg9NwVcSH2SsQ6Bq7GQr5HTMdgUMpiT3UYS71/HpfaEf3xhz8
G1ZaBMscoMqvrr5zgrGy9jb81KD+MMYYMA2S8N0v8mBpykA1w+cPuUFHZNPnBax3
fhLTkgBfPQRJhkBQdjgV5cB63Cs7Ba0etCVLWbVvxyYfV/Ddzt0skOTamFiwBVXd
60CP/EJwcsJrXVQ81r8ITqkKnTr1n5GVQ/x0koLT2NZxw9PsTeFjZiLm6HmCPURP
PcPzpCduS+pYCmIXn8GXOzaq/59/z3qtI2Gq3jM99VKy4lNCIaqkDwdaDtJCIZ74
KlLBdfh5Scz++jQPoX2ObWBa5vKhYzGzOUlApzVTy+Wb05ItXrD7LoWvy310pCCe
IFrngJEbyh1fCZXAADBe63LkL84JJNHrL0Qx5KHRyRSa1UvYKZLE5edcZs5hSeCs
dpFrO4S0y9+KaLXhSuNT2ebuwi37Y1qnpXGTBeGjTf9sd1dLllHOBlzMVPzj4cSF
fsbiIGntXDb4+Caqd/oFNgXPG5+2CfVJv1bJjZAs2ZapX4m9s1vQVcUmJ0d7JO8h
DDLRvilOjMM16SR0aBB3Sm/ABydux0GlA0SpBADkFJ8fujHcee8ACwTM5aQVyoV0
uIEcu5Nc9kpbEzOAtbOEDM715QcIJH7qZXUofX2Wxn+hOGf4lWYtiXW0ikHmso3s
kZnrlX1uMMYoWcfzhWWl23Jcg4PeW8wds5jnIVkFS2F5odC5wKwgh4OoLz77mm8l
Ot/LUJcXOqG1I363bAsy8KaAVeNiulr8De3HGN5D+LvUyL51YkTdeINRBKCTYiI3
aukYNCILxRWxCxoRGCtK95tnegxuYfAEpmMoxuTUKr57xap6z/hV1Ugz99127PZ0
J6S4UXMhls3H94ylzQpijQ56MiUUe6EgKRAXHFmKHYOjgXCPrQh4KBk//Q0TOhSj
pNW3Rau/q3qF84f/tYVMupFJXLsYQbd1PeToQ19GFU8w1M7BzTV2Q5iEOVpw0FTc
m14HGLlxGgS4kvrNcp61SS8Y194JpdifCT0CIH0qi7VwRGIneJtET4yM9H/bvv/L
mGEHxuV5CNnuLEGWgPv4FgiecpnJV1S0erXMu7x20nrWK4nsnE8Wvvcc00OJBjm6
VVi8CYUsS688e38WJJ59OG9FnlFuGuNcvCqGLwmMxKXjJwoMxFwjG+hr59E26Eq6
EO/is6q4YuLI8HfgDkKAfPdDyibw1AczPV+8Ow4ZaDrcU3ZrzuQEfmvOEir2MJdE
ib4aItqJJnugHCLnVA/t9Ggls1Lz7yvCn1Xg4Hh3O0flHwkIAuYnebxvmIQY9QFJ
Su4CQU6kKkKfrrz3r8y0v6jyNujU1n+dPfMPk4cZ65pw3ugptRjf4srWIC7rBp75
OVX+z+TdN/wPHM3XCDJTIT7iTHDj2i8YTDGwGcs8XUs0JKtRcudjb1yCmp9w5Ijk
FquB9AOni7fL7t7cwdPD7PCiSmzTjd8FcX2hRZmwA85w1yei1+cTvHb6KeenyzqF
6ze9MICpnqpy4CPqGwDAQMhinwYmhuE+GilVj7GDg12qv/uzZ/cQzXzo6vGTOYoG
CrFdf5OCF4+erR9bUlW4+CN2QG0m+og2/rhYaqTK4iHLnDmtx8drAKjCjJ5dXweG
1zIblB1Hh3Y/lzWPJLF8MBJQeVbuS/wedrWuawYD5rNzMi3AuRsNv1ZFmFFIyyDX
HdZEYmOQrSneo0vDJUPeBDdUyLl4EBoj9Bhp88Oh4bdJaILjyoNgjCj+5vCGCoE/
MJ+feCE0JVWzwKz8ttyArTnHq2Ks6wY/CGebTBgH3M6YvUJWwqZLDsP2Z6XzqOoq
D7M2/bo8O46g8Oyyw6Fw1Tvy2SMtyzEvm8uqEURReCPRIew07CSoq2l1j9iPJgYR
PdFIhg8HqEfElB+1/Qa6y27GocmmZPUOUgu0K9fHTH2cAIjonasNs5xRbYMNZVHS
vTeMTepDWfU2y9mWohhzKqi///kfWaryJGEF64zjM2IVI6cJbT13Vchd95D7J0eL
M2LLULpH2SF3qWg9xuMNaFKOMrOcoHD5BdBNKqNhfq8MbuhS9Q+8hGskk87t8SkM
Kx3SldQZBFQ4JQ8RYX/1FUd/TYOZ1hZI1f0yMwWfmCeE9Slz+E49BxBY/HxXxSTA
4Q5rGhJJf8hVLa8gw/Jd5V1d29sZpPv+mD9v1OUYgqohkLde+8YY9ougNViL/Swv
KuxUGCQKgZph/PBWXKahL7oAkAITHWGYVvIiFkOr5i4n+Snsks8lhwpTgDODNYA7
IxBWYO0517HXVv12LPsqWJ6zjoDsAlbYdsdKHXCCtbqY5KKxhQDFHjZzv836W+TZ
NcC9F+EIYBpjUhn9R9PbTrSd2ELPvuEfFYrALnWACjkDeM41txVZi40QLvZ0xv30
fV/lIQVInheYW1DLklQyX5eiDvrzIQGbZhgTfw2YSraGwbEsUt9d9DDXFdscNTvZ
8tLJIDfhJlhl/mNmEMGylJFI4Af7oXXEKkRpHDxlsy+Dk0VFAybHcJZ9U92SvTwU
+XbNqkwHC6O0dvnwB2VKk1iAI+1ZwYQ0WBrxGdgiJGog4UP/niav8ITqi0eUgDX2
oz26JN6QAhO57//c8zu1yCkSxhatZLwUI59xaYahFeGFb9Yt892tv3VwDbSo7hXT
mt7QQH+CFZEyeBM+chS7Ggy1crw20FardRVz5zFDhf1OhJLLLTyVFmrbP7jMDsvw
k+VhGaiQGMtXIZOMOr0wLrBo5qPuVqB2XP2AgUmfmgN0njl6Hj+Out1omMyHy3TK
g0FgldveHDqm4LRs23wuJrAOWazPguQDUJNwsfw4I6eKU2I6+m76GLX5woug1NKw
h7J6Z9cCWDEQUsKDTnoRWtYDBGYuAXR8AhLlB4L3bn6vbPOcaSev8AVnkQtCWuqQ
FalhEM8f2LM6B/FHLpDHw4wl5uGLbuFtDe7w1427EutJpMgsvEYYclj28mnTrv8I
Mtw+RPATrkgERURHUr/Q+8ETdF+w8V1FrwUKFDdDnXj+a9T5rHjKYexj8YAgPLqu
tPWqAwvN87a+gZ6vLegdi6izgFmDzoUvJQnh4fOFpxSPNYFmq+am6oQXnnOeoIY2
4DEwZThUbjEHSHxXFQziiYFJLEjuhjaB2FBWLpUv1pyFl590YGsETNc4C2YLM90C
ly1PiYUNP2reeNSis8MOJm5V7V5pIyga4gbQWKSRwfBftPgIvpnmdV2H00LQa5OJ
Q5Jw3DXMHilvJ0SsE5I44aph9HVnUrwn9wF4kZMjsM73vHaIa6mexaI/RaauqCgk
9sA8fRGox/xI0/WOVlwt0eUwUAcuRPbst6IAzShTFmStjDzqORLpyh/NHXiLasSm
Mcv4GomsQYeVkfAv0VrtMOb58TQs0V/liulsa/rKrhRBEVxewxy+wJ/uK0lwuUpt
FcM7di6Z612sxLVeaj1j1woJzS7GhP3X40N9Lwdsd452ameIF9ioHc3JbQbHiUjq
VQX88b7DPevTuEHn4Ne/ROR3ek4O3DqX2DzblKK4nB07/Os/dW4AkNto6NDEvl5G
fxwNhA4RqpoOcdoeNBDrszziumajRkH+fjscl7oK00s5jf4c1AJpi351JyskNXw/
5N+5uXqXFIXk2+tmKkIIsesUs33s7w2CKD3zcgec2UzzMV66HOhHIBCurg3aoWA2
zrimZRgYI/tRGh4lCPhTjNVs44aiEmP1CcMozKx+L6tzfeIDhUEodwmYtWHB9PsS
RDGxCgSimHUXjR6qre+vx7XeAGVf29z1dBryfYMggecGSC8uWPE2naeaxMZLRYh5
XkfckMzphinIG/u50KHoJGvqNkzEX5LMl5KU+eCALsAHHrzolyyxxATZ+IcGJog+
h/pSpXeeFaNrm3yLx4u/rBdm/m7745wKlx4eNF1MpNRGXthJwCjCNKF8JhyL1+FR
JToxgwZUL+NqE01R1tTxBzM0eltNCj01e22ht/vP/dBsU8lgG3n1vbSlnrKscqYt
Kd4TVqWD4GcldeA+M+RlebBMFC9M8um9EfTWTukRgGWZkR2IDeY5Q4AjpXvG4nCI
pamOqh4JNCqYIz1dtYn27UcHjm2ARmn+4gQxsUnKd+8igpu/bhPArj76oFVV76Ue
cSrCV1pfAS87X6d4rExvMJo0Y16pOmmt4GVGQnTDhyZ0CMVCxjTttoklEMDOZef7
koKw5UG1obzsbVP9+vEUxiyS1Uu0JEq1OlafeA+LAxalIZI2rp2n8JehSc2xiC40
5VNXUfbFSQvN38YMOI9zsgxSkkxLt8wJ6DS4UIWSI73iXBkft+4GMQgMy8LFAaCn
VGE0dNNlR7qNKe1POhHL9up/3EYx3V1axQS1vW8yngrgxXJIwJTwI/PSNws9GT3X
4fyLrJQ9qeUPYvRk7eNIdfufxTO4/M6ZzKAULUj96xeHj21G1uxw3R8lDeiBwJqR
ONY9w1rPdGQi1lMz/rHxt0LZ3Tb8d5QY5ELNwuHb3Fz3hr9U+fne/RizvfLSxb6d
zDFBsCHNxRHaqWBDAMNK6QnWViTf1kKvMAqppeWK2T86t1F/JNaPaq2GVrAaOCpy
VGFYuMCsK+Av24TIDusj1FhmBUp5TGUpO+SZ8RyO7fK3HoLH8ryWRanOLUGm1W2J
No4PmGWcKa8h3sSIgepzwRf2eifV21P293QamhpW1h5EV52G0uJflEQayE6Tz2GS
4hBlI5hbB6GEDq8qo1VrGWFmFcAIW+Xvr64/FiMqrEaq95Uzj+UGqR/NVbo+GR3x
dqs0Zb04YBTCawA4Qa38YHZqExWQtWufY3jXdW3mrKmmMfnRa+TE63eTEVVvzy3V
lo8MXxZSLracBq/ryXK3AHNwGdWp1+M4frjcEgdFAiub5aAsSEmjxp821+k/whtu
3pX2lfoMpjvm4k++p+mXxtJ31babd9d6DXmBGSEMAvfFSjPJUeXNVRl/bzORwGoE
xWFmtY1qkafJwBpwYG/KX6BS9QYw9UX+0XmXtl5ZEeB71M7nphBSyUVKc65Ms0hS
MdwQcA8xNrADfZbgDw2TCTVW+45pX50b5lJcZ0Rua475Dpnlm4woly04CTKrVYOe
R9G7fJTSNIWqkUNcR11yS1g4IPhyDwzmLu05wIohP5K8Eqmw7mYpTpdeCfjx/+ok
ig3I3vOv5SIsoJPoCO/ujFRe+m9dUTiQkcoIBEbXIQokiKJ7yAT+PKWMkK/1VJvj
1edqBROVajQhGgf5yvw3E6DVTpCGQ5/KDjPk1iO5IsqRbLtmmtGa+L3qHBXn1Csi
CILaAbESkphrCQXQ25voAZjqEL47GTGfuZQilgI3hZTN1xoJzJ9IZ24WOz7JwWEQ
XMiohWOXc4+JM/BwCFjZizAruELSyNgQbuW6nScCVnoFIUKzDQzqnHSFIvBmDiEv
6MXSHMIyh5hE8F9PNMu48VIZXbOw6YBm3cq+ZkXHc0ttd6VSyf0dQjB6Mei6chmv
GSg8gm8s0VPTua42C0La3k80I/ApeyqgzuqCvyQz482ioJFHV1Wa8K8vlH2RHZPj
SmnHYmXzeNMOVIl31rgIXh9v6uRV/xJveGZcZ475sgkYQEozeoA1XDHIP6wREEmc
KY5NOsJH29YMQnIBkcOWzeSXLcKLlEpWvD9g2+iPMtPKwajKZg1BANKD4dWJOUKE
kPuRjlyvV4LYww3mMci+gbNedKODVosAWLHUpQMPnyPLPMKBVxA+3vCnkej7mCgf
V/CBZj5EHT7/tUV6TXw/XR1fvEe+eOPtTRMUxymEkH7mYcoCaDzaiRZqZgtoW8LE
S89EvaMTegmE0KdYSu8iK8WreY93MtuwvjdY61I85BRMM5FglvfYx4YtxdP1DVRd
cQfQL/h5lzZV9slD83iLKLk7Tl6rBcojJYsclCzj8ExiZgYi9Bfls0frE4cVBugH
+75BOagPGkq2hth+/l092phzTTFe/mAGDMyzoOaoqfa26f8y7+jRKH0/Suwf+B7q
QhYEKdyLR4m62fTVfd3RWV9d6/cB4yy0i/XhppS6866jcMuYcRjtJOh8MwapzzvX
OlSPcbDkJ2O66V63xx4fw9+DLmUtKUYRJb8WsywH9v2rdP9fKRqTEwqclNV5lxgf
k2rGbyJ3qjrw3skOSZaroXggI64TfN+i+tsXNGOF9Yp1sAIGhMkeUEIMBY29hZQm
V0eWtopoOIg2KRRaAYM8LAWVLEcyH+IKyyCFgFTZbeguTQ3zkNPGPsMfmi20IT+e
wLhOeExKH7RXtgdTxYV0ms68DkRkSa8DslIrO45aaoAfkO8Tl0XVp0Cd+7yVPYh5
V00n2Rl21VWWB/SpfT4aaMr/aEmZtFIjn94bADLONU44JyLy6mkvqRJDteiyfCaa
aSpHL6SH9v68S6No1je8cCj0Wlrer0DoFLkmuOOIqMV63hcR8L8rX/TuEcOOa6Ps
xx68RXEkE3j3MCWyHgdGUhQasePGKT6JmP3UCRKkMCgTPjJouaL7c6brnvcTRiEI
k/qG8rAxFg/vmBMvR4wGjE6XUswX+qe0lXwzVb/NLZrUOHqDlPwEnCWdgPALyy+4
4rIOfKg+EZfUcitz4En5aqVNnK8SP0YrF35uk4Ohz6AfsLlRXAcnxXgFOM9ZBJOl
+zvvm93fzbaheuf/srSLuFmlAJJzcO9pGJZo5SUs0DhkoRuEPJ2fPEylJ4GQ4oUE
Ltl0fU+4elZAMzb7f775FLM7fEV9u0+txsTG4EwDcBn15q80GdDr6iWj/QlcLdim
hUbBMZafH32emPVmivccHimLY097LO7AFBuPaF2X0UdRvV01jYYTIC/fV+ereh/X
o3xKtWSdTU5568/UXf41QnIChDHDolnR8mXNqNAx1ZlCl/QevuFGyh6fa9V9kII0
9VGrBxHuJw6STJZySj8nVXo9AKKtuHGuVSe5d0F/xrZ+N4YeZnDTcm+drsx52oWU
zrzfDFJTlE8H670QLzXsgjueL51wyTNqfuVKkbMtUCGysK0K4+lygVdVw5Hn8CBB
bw17QFdwnHfnMO88gAoA3oLJ0LmH/IoGy/Gvz0PAHroZcdYPWeuDh5CGSs9YoXvG
syktQsW3/H8V17iU50UZ4RgHXmsEc8Ks53jGKHoEaoI88JnSw1FGkHzlBsTTrMQG
/Ybleanxqn5KSUnyVE9jS1C8gKIFrw8J41iv9od3f7ogrRswKBKujdKWjV2zuPcA
0e8YRGjeGBDrlseUtGDdMN/RRpw+cql1JXmp9iTKj/Zk6LzzabMTnJdOwYvXS4wi
ptmCOz4mo1PtFWQ3XE9pgschFdrtx3yXci8n8Amuk1EcJvtShsxC6pvkvS9lb/Ff
6ZrTwzAlYCHJvDZEu1rL1x5OV4mJq6adM+5cHmYWgKywXBPmEDxQnNhfyet+YJME
CEJvASsPGdMGcLPFkAsxHp+uDwsHwm3lEEUDteGSng41bEh6YjAkzIhkMUV/kOY9
tO/uac1ggw3rt0xjQL4z0RLoqu6mrJYlC618FxqVjB0zKSTYkC35FzO8k0i+FNuk
WeZIO2qNmeKEH76v7wSwXCxUSEPngroYoVKcvFFohWRA0FYuxdMSpttHFPe7LM/9
vDE+Hm5OYgsaWW5KtTmiquV6dtJUigXsBF6dgjycbkh2RU15VJoiuwnaU9ZrXU6U
8EpTkjDwK3v2CNpKpraRCcHTvcjizFyLVIRU+Uw82c/nyi0i52r5kiUWGRpS5ozm
oie5Lrco6SP+VjrTxj6o20MqLm1ARX7mqk2eA65jU35sDuySn+h6fW8/myEQJpqV
A1L0fLNmRB1THYQanBcEqSHbqhqy6c3TpEI4DjRclWv0szv4ZkAfYaSn8bqIFHuP
bBmnuAOw7ZM5Q3g+966tKTAkzuzAzMKw8WF/chf8FkzY6gJNyZnQW9bHIdTzWspo
CK50bHhUcYn0beapeij3r3lNP6jCzmn/xdR63thc7EEMZ4WIQ0pSG5y2/QFfGAZ7
t4ae1rLM5/K01CUuM8A+z+vbq/IF2sSZA9na1N5DaHx8sjGPGWZePXZ9oGYxdGSB
UEoyb1qbJae+/e7DUUdNyEf8MdvhdoDmdyacjn3W1GnOd/Tq/hlKcwmC4hUpKMgd
eGxuvfmcko44KSBehBu1czJk8A1CNbwVi+tGljKOz+D74VZvpkzfu+tG2qMW2Zk3
yo94FsoAeIwOy1ppA/VNbMUVz8VxvUwviDOeqRGewQLeXlrt9gZAwGASVVn0lAIu
llUU113Du0ZtBLwLx5Dk9ad469UUqyrgipuezdhkJx5xK2veTK1a54xdc2hbkYSn
HvRZH6aIhje/i9BM/YtEnp51Gl+oCDbR6O2jNx7XAHtlcYQbPDBxSsqktOFVHgEy
5WF3UbejuAxSwoyu9Ih58HMVO3a9iSty6RBqV9TSNqQhqbWn8xJRtOdgvWgHvNGu
DyNCD3YbAej7evPtsq1aJH6xBm3U6Y4nlVpn683V1Y3IvALAZC31kiiOUGKetSJ0
ZwXPDCwl56fzFHFtqCg2/vCN97NZt29nivmCRuSCwglEAxqrvlCHS6VTgzU0OF40
qMV5h6lDAtgaJIf3BPe/ROFbSbycr93tk6I25flcCCO6Ey1FGvzHHVWO6jKUkIKi
KWoe+pnHmH3VwTpH5hiXI+2Uf3UDkW6zPIA/NTTg3+gZnL4rnvyNAMDePz9gzP6/
QQYDabaLOZ5Cugx7CIEi/fzr2GzT0+Na0YgE0OvPYWhZD9BjhO+4FDV9D+cOJBpy
Iip4yAq4h5BPldsfX3lCPP6+z3Z0ojRwe9/2CKcjssucljqFCXm8rvx6zc61sNqn
ysjRe7tqrUg0kygjCBKBe4INYSOIteAaeDzJmvf575MVF7OiJD18AshB+IMUEQN3
aapCncCq72Gxb3kQEhcbUB6L7D0crKbVn96d272g9O5fI5hLDKhxX6CcLskb7Chv
TGqFQrQLgFZRxt82ezar4brHyxTUlXXWxW3vnkympKMenBTm5Aj3pLm+2qi+3sHj
NZ4JrWVgrDMMoGeLcKH91W5jatQeprJ/B/pZ6g3h5r/ApZ5LlSMoR5y7RA3UQo1r
i8irWxrOMxvUB6JDhGBjDfD5YzpfzDa7KCOzh+ozFWZNpjgc0oyDbxwmkjL7U4v1
AJApWZVAHEDyIQEjs+GFLB/NIGCWb3ZJLOm7zwbAI3A1vJ9R86M0Wr7q5ia+Af42
x3E+kZ5I/p+aCV+9el2fN2C5NYZWa2Kf75Sxji4cmdq9tcjE9k3KuGASciQ3kqiP
JFWpKoxU+QiB5NEXX+E5uzFBjTV0n7U3L0Lymgt5cT654hKx+U9IUttzgEMZoPKi
b5vLbqd1M5pXdi2bfaAoIuIIbiq9c0loLW9/KUIkWFVPMoGxmsS2pwUQi+gtAZ2h
8zbt/zwIgzkfjrq5AJ2F7GUSHyfraQF8SLT9Ct9FFybvjOjxiYtsCMLOVnZwhe4Z
uTeQliuYI+9UsGIS67sq17hcqOJFQ1V7CDNiOAtr8l6HpvlCTS2QMTXcZgLHOMIf
r19FrFKlmbfmGaqARpTBCIBe7Av0EpU7nLsZ4I97wEISEip7mMb0nEm/5orea3x5
mOeutqG3ZM0E1i5cyUDnzsdt++Dr01iC6F7/T2lowR+PWv0+M8paAzT5R3ASX3ML
7Px5BkkQHUWJXuDhtyMgMUEuuk1ecwrzROgwz786kR4+YzCT8Z0uiYQmthnsVSFk
Zt8lcVPNgoXafjPGCxiEGY5GfOAnD6v1mnAY/ODAPZJyY3jRTjxOG4Ki0sNgcEBP
xmVMeaxC98qQNGWJa9Ir5HKF40scbt6HcjrlAw2RaUr69PtAdXIf6l3pehfl6lpL
7xpfF/T/v5GDxveXY04vOsBbO5cKFdbegNfCE6KpZR4a1QhSYZfMx/gsBMpcC3mp
SimGqzOOkxaxA0IObcAsCYZsql8vNj5PQHR/KOsYb4guPwrXdH5MtDHM4PjPXjPt
ktcMfps2I4FTJL3Cgd6xafNSz1hOSi0iO15vUepCrmferiqnvGu8SbvZPTRGD74I
lAi9Z5bH26Kt2lyTF4IEkFbc+ER6VJzR75m+/C+FfDBlneQR6FE1/fUftnNjpoX0
MJNxrwDRaCn4bQqq3TnSy6OjzHXCKGGjgY44kBoHiX1VRw8tbU6WfIHMUnQ3n5tw
KpNZyWPLQ3dHsbWLcZO8cTIQqqA5oDyrmncLgLv06oZDtnTL105JNqXTc/vAtzLc
wq9cLwYrc09vb2+KvtLCmRA9gh+isu7JH+FrE+9zIGX8jS58UsWIDVykgiTIlMC8
KmLl79mJdoiwUHcRlwOaKd7kZr0hOHvfDOnS8G0sjEed3eDMpP5Qaaihw2NMTBqo
kNrPt2MyfW97emHfp80DNf42GfjGWantBdy9n7m3k5ZD+PTKU9xypx1TtT1atCp8
waAPsaZWrd3hsMSXvTUMRXNjP5l5DnIrkfDK0Wanv+I0YZN8FTCr9AppRkACITh5
YaIFnUwsV75+mOGE4upzC+XzfIWCS9e7W7EsDnpAGxZHpCjEvktV2zBHxcIkMtfu
fn5yc3nf5NdQ9TPdf1bmLXUwJkvcuzlWvjHY+C3uOwBPPQPO9v2KoGHGs5uug2b5
LeKT3FcSGP2GU5bkbfNUtj2hSliuxdpkUPGqj1hOef8wF+9BYLTaRLnVOWUZrvEV
gTqwOaQsjAjprcj9gEHV2WwOLDuol9RksPxBSS9eqQMHZmKDHLBRcF0C5emiRbRF
yydFQlJRinMJN+Sevhs1gTgKV23M6PNqJyU1AH8eu+XHt5ju5ftrfSOHuw0b4peB
z/kix8iEoTEWel2cWf+TPrpThBXaNkYpuF/0P83iTaeByV4hH98I4n402Nky/q/w
AdZsXLLJIy5ZQEAe4sEOni9NVAn90/JsTwyovpSBLiV5rStbeuPFA1VYzSFrq55A
yElH7NxW/x3sh36z6ir4JllLLfIWOeoZ8Xm/fwrYOk6Smd9++G5hGAktES/zRLdn
tSvYthIeN928FT08l1BHgVe+iu1KtWMqiNpnB9yikzjWHuSQdhMHW6K0FVww6diH
j/VZr09uGdLU8TZoYiQYC27wnyzSgs5jpcATfrPanBkWe+nnVrHA5wsQ/JUvBGXl
piyUVU1iwvzraV4XuEf0XZvV5mo+7c/WIyk8jJUgiclmQ5Ti3tZLVcR3tjJEznWv
neqdQCT7ZCX9VXyXwRb/H237qWrx77EBj//TITKh97P41BLELgoGP07ZIfZV2vOx
hV8sCrNeQMu3NAFclO7hreg/zntTi5Gx39+lxi2OWBL8Fkkwbs05RHS55So0I9jy
Q3HXIYPvQpfhCjqS3HqDWfd6qCmTjLtjJGs8jF9KQW3LQPc6v8YbBiwstPuA+bSE
3H6P6Xs52yZXHN2x5IbszFbhE144H+ypE2Z86l8SsZiGMiLyNNIBqaojHUpfL846
Ap72I8Ktlb2gJEiQx8aRQRItFvGpg1Wk/FT4I0eMqe5GyyOON2R9AVW/CvntWa11
G8NM0eBzsnrk3TDuwbYSJVBbKQd2Aq4+NVGKxQASPTzcKp21PCBEBrdKOvd8mmX8
u2ODVUIS8TAe79OBWsoGtMHZU9hUTCeAoWrULLbXvTm3X2ZCT1wUIrizbE6fHpMY
Iv24IGpO7njlrmr9+r0FrlViVq8ppRv3gQ28apqthzigDeseyLoh2ujAwngcjoa6
7pn67BngY3lkdjNKvcxX12cIcCpnWU0k6NooKxRAccaShMySsDFzs18KXUmj4RTR
/1P7gXCDo1BtECYfyYN3h3l/ySxAIWnmZn+TXV4efcD2AWFmKQMyXX2xt38B5D6C
JMRp374OHXaUaHn8Ji2yoY3ONpwKE4WD80m0lGGQV5tk3aIBDf6qRVwCAkefLEn8
xnh8jHEetycot0A+DNXN/xgv2oLo3KQ0fegCYKKpCwoMVZ8490cGRBP0zaixkuoI
Fttn9gMM5wHFN0TI+NEwTe5yh/nJ+3D+y7rWGg3GpyXxP6N1liTbP6TbuIWhF9Gp
ImSiVvuq/Q74cezVMQoX4mtGS979AisbLn+VBWkpVIwr+YCl9IOc8jjwTi8U42Fc
m1nLkvd1QeZhQVq1R64EqOPo7ahPpYrilr+xBgZ1Fo20SO9vksUPFdTIdSPMbLOb
jK6hIGBiUE7X8vnxtWKfHh5I/oPH8EOefj8dXpE+oQeZiejTAWFEGzwapvxAyOrp
SmGepS+B+fZGBDQqltEHwQ7Ojj13EJji+LCSAdDzhZM1MxwJmXAHmJr7l3eSdWA+
NlVBjVnh9M/2hqgMiBRDO3rXDpZ6ozUCl9g0MxG6THUbM9BELGJbHI4FUMpe3to5
9NBtdQ1z8nQjXc7DRBkVkgH8bqk09g0ZmyoKT0VAZgwLJ31uP4chb4ZWTuPj57Xs
9BEn4a5hyYExVIX0mMIOfiZ4YQgrT/Y2ex2Bx5om6BZHM5UlIh39LO+OiHO82trK
WiYsKippnXmIl/4tfExHq0STFIb38MATnFIT798ddNO3+nE8jMi1dVUXfus5n+4Q
MwzT0W0fvaPMRy4J7Gsor6hhkVHJ436ES+tjk9tyT/X9P2hYMHqflqwDs0gLiR0S
c22i4kCRX/Aa7pXMat0kV/D9v2nRQcjPYKwYve0GLVKWUdrHSiRw3NZCm8SOQOfy
6Umr6Lez7pqIHOfdSe3PQIVOFhPfIZzNJNUeODEZlQY3RMSDpnOWdV0PpVY9r43T
d7Tefa3f+a1l/ZIpltbn11s7uNDjZBrlRrzhbsvwIN4TgSFpbK30yQalhAkVwJ1i
0xR48RFV9ZyuOJazHlUjIcL2ssvuXV7Mc3ZBkWLopdVVocOAnUfsLjZiffIE1IPc
8YXj1CLItgFXnPXHguo6gDdRJ2McBrMqDD68ri2Ug6Dki0V0nI8dKIhPpq3GPIfF
1UZMLMn92TECYr8LgQhl3Q4MV7KkWzZYWRVqgtlNDhf96YxFh0egVAj5neHBQddd
trDImwBRaZ+0O6X6E1tuM3aMUt1MG1Zs/QD0isxhuQrWDSnwBtGGNWST3NzAYVkN
ZZ+JYTSTSo3udFrsb5w+zXyqcKLbXWnJItDV8axdmqmWgEhDRw5kKFH/f7fanhm9
ze1yNoPUoJOd5XKfjAaKsccoCiyx/RzSuG/fnrAqadNkREwUBoXfIXnxbPoTpti9
nby20a6PkseAVGAqBG+2LQQ9j1mmXGzb/Bzz/EKFm4CfwBMW97drv4RFC2s7LDXj
gVT520ye1DHpcq462GhkOARQnk/1mnxw5fhbU2x/XvYNgzSOU6v1vcwlCLqI/WiK
gtk4/MhkGGxYJaHnJzVURMz7Zez5kt7TTAP2FCRZvsFCrLlViqy3eeDaD+zGMoP3
+lBiMxO4ZGDAqP9pg+7WOscQm5pDaHIipFugYn9t7Xkql64k2WGHLl//AM8UgUt7
cvfGJMIJjMre6HrFAMv+cU6K3NkfXhJUQZkn/LAkiUDuqM0mnloFk2CWgFOwDBF0
U3D6bcTfOptkhS1Gt4Z54fB0TeD548jD4qu6O8AlAyJjIHl2WTLlEWAySTA3R54y
T778+bl2YpgaaYqMfozwCObHf0SkhvpDV2+jsKYo4lwanTzVk6TslBqI6orrCiAZ
hN9somyZosuBh0sDTC/AiHuFKU/mK1JuOYhLtCZ4EmD1w+c7AdL1mpwD2VDud1Ws
NjJNdiWKOA4iKM4Q6/bn8vSbHh5cTpV90keeAF0yNA6e4PNFIx5BMlZ84AytX/x6
DoV4ljJpW1pQOo5hUdXgTKcleEZe4Ar74RgxT8Li8PDnz45NPjgnk+w0rB6FHiGZ
qzVK53mYFFYBlTlR2MZEIbC0ECHBXOb/TBIy3geB8cEJIvBXtwmrlFahn3SY/MGI
+CF3+qEsRKq3asqLRm2i+UO75gISUPHWS31JYlMtEIAxdAlKpiNSk2y0Fx9qMImC
rtY01p6+NYYKJG8ykyDW12R5PC9FFbV1Lfx3HNaxHTp4wkX8HUk2lI3rKX3R5XcQ
mWZdS285lYo+RV15WtWzU3Po86Kweupkpgb2yjb/zjLdr8quAjIrtGN9ev682fjK
xRWRyzIx9iepsokT+TIvNONLuR7uYy2QOzK5U2su90VAVT04zWjM6bvINIIhpIte
U508IIkKyFk4ST791sMuFf0wAP1SygleH0e2rDpsNqMdS5dBRhanScSaYpoUHV5z
X7hGDsqHBRXhD3TQ2ucPBgxCV8+hS+G4biyPqEx6/MPaL/dvv31B4X72JhukNWmN
CHnZg55R0V+UM9c2Ydd4/Ns9nu/hP0LHTLXMaJN7Owb+bZs7IxZRQoBv58HG3USM
D1gz/7n2wPgEZOsOcK5C7sMmj5U+oiUvYrpOVsc7ehNMV1D+jeZH00eRAiq82BI+
ti29yukFwi92Okuk/O1BBRGt2VWul4rpcjztPnYEyzG0Bqyw660pFfH9lxc2YdvO
gR6QlOYipNPyoYcRkEnIPfjG0eQrlT1MZD08xxJmZ6UByU9jT5RFfKn1rf+QFJmB
TyQYU2houHSiP1ocxTtKlUW0/IQZEeqq/zvlfivIJXjh+DCSvHAKZjMYNiFdrBWy
CvkE+nxAB3eGRh93x0q2t43sEuL5v+8uLrcNEjOulI6edLXY/kTooJN7UiZuF/Yt
x5UV6mPn9mxlk8Q3o5tJSv7mhMUQa0Ik7Z8WwVaWC7Nfs3lOtz7ydGf3+u+5Bioh
2SSLOUUsmPataXStxJtzwvdz5TGZXyadwC9mn2W79DVbaO5OP4VyHHJQ2ED2F/Zj
CwzW4fcsqgIC0SsU1US8EDPj8AP+msUzyg1dI51/SGK7XnGoVt7YfP71at5C3Gxh
bsJ4YpA7FEuxzWZ7PYQAKnuQVChV/VzoNtOuVX4Rpev+YJae4AGxyometF8DhOmn
SFxtu2LLa7bKU4m8D9cIwqFyyWTd+3FhdaA9ngbNtlCteHmilzzsSP6w7uyr8rwv
PCNS3OiuTJ8UaLtDWafgnIahQA5GJRaR+fDP6E8Uf2abe/4MnWgnmHgKL0r5aAXe
2oM14Ock+bKA/9N74MKXYahzASOJMCvPYuk2r7sfRHgn2ZGhm2/V2bSNRYXZsvMx
iPl0DzelrvFyxHK/qO75QbAhtF2ManhgF8FlK6VuxbMwvqKqqi+TBSWZuk67yBlN
0LJtma9dLxZj2ZKPKLk0eNcpMraj29Uox46Jfkcl555o6CWF/T6DIPIEpr4VsLaP
cMXpE1UXJ7JftkjruTcnLG5CzZt7wQlYI6lPjH/0mqwEZz/aWNh5TTsz4S7FstvJ
KJVeM7HMdNtL78q9rt9/5KuqeJsnR+obFhKgcjK5+XvPARVlcFAgvUu+mvKsEaU5
7ZNmXiFW+6dA4Zlr7z0z3EKKfWC/et+5PGHqPgaW16OUlahOY1UjB3UCeYv/piyM
oHHvMuQhG6fdtXG2SfgG7pHiD9Ihd/d/OubfZyjIpp1ouD3K9k0DrMRs8qzP9K5N
srQgUvtbvrLn39V0bX27SdRlfKb4xRrabFdM1ioqFbTlZ9n+k4AIcE+R0oRAHVMY
RrRqvcJo4ZkipMqO+oJ/LbnLoGtnrtubEyrlwCQ4lslqHgxfkbM5O3YsmXYYbcyD
GQ6xowGT3IVMqHtMY7h7yR0ReR7vO2VQRr/K/3Ar7HsOVbzq43cv7VirPjhN2A/1
HYKQbvqaIlKkIBiOoBBe8Zyz4XxLNciG+QhzmUiyD1O6J7MdRkHLGxPO4t1ULKDF
E+jXQ3rCrMd5pzosMMFH7MYM6bmIz1C1bRBFsv6GZXLVjnMm7GFXLN+kwNMS5/cZ
kO6R9UoEZgA5zmvFmWqv5FU6VN6CsK4T73YvxfEqIuHfCXv84phJpeTXv3DBmhZ/
Nd5i3K+fXtqaZo9b29KWTQrdRijapfgU0zTrPDuGf6cy1SzT431baUINM8uHspGO
zWH/9pnSLZtf8JR1WyykAJAFKryBES+G5011owp9bR/9OnEOkoxH2fYr1nyvCm1L
i5ViVZnErs+46nEskjrva3yy0s/IuuLxcDMVzDHr8qCSL1UBIQWkTTJ0mPo+meCo
8+lzK10+PCHvMuZF2TOFxXLgmxygO6LXW1Ma2K1Aurw8SoLED3x7lBJhfdGeJFB+
jfzf5Tvai/HBlH0OJlx/nWZq1BlsrTMKkheXGj2kSCLYdhHnYHXiIT3OmCMTmhb3
mh0+PPSxQYoTJjKyKi17L4H+pCZAhQb3Dn1PqUbqUvzazk7az4BatUo+vjQpwJ1A
mQvjPUVGBhNJzy8ZZOaBiwxTMIiJ8bv1PQe7ob30vMRQrFdo4BCefyPc33epsxuv
ikdqmUL19A9RuIz+rodR0PGFug/RWGQsOn0KP5TYyp6BZ54HJFmwJ57AiU4KHBL9
SUracAvcu+M5JKeutqdhAu4MgcOD0pDudQZPEmZ53H96biq7k3IyuVeUnFrY5QZT
znW9op2H1yu60TCRWsE22p4veHhbOMfizsaY8yPhLL19pmz5LMgL9YV7zVAdUIzX
KR0DpMWSw0zTZUTjn/gP9b/yBjr+p5ljKMCA1ddbFxrFkXmp/P+UHq+y/foS0hM5
sY3lTzx9zmuUe5D3XViest3GpV6SnUUdkQGgn2wJsomxYuhnORVcsOLFVwi1TClQ
T0+fuXdkmyqJgN6wB8jnxsevgBOzNdECdwgx3liDCrx8MTdKAQIjFvhOY4d9cHT5
FXh9WxX6Z2tTHFTkU1cQgrgtmD2GdeMJh5qIFj48aAhqEF1G24/xQCDo9yw81Vp9
PPrAiryT36WIVmtc5n6CYpmQpkmBVN/zXamJ7Nkf+jjv0b2p8O2MwIQWPIYGk0Qu
5zdjGbYkdUgSBB17/PeQU0ZEaPr1ii4uJ6oDZ4viC+w9nbLcl8FhubPa7NEhuynR
R4qfkZWjqkG2CzLGelUip8lAxxu4QWKOrJjiIJ0RUXi4LU66ThI0Z0gSYSwPMMlT
UyZEWmOLHGAvtqmREfuCYNeqBUX3MLSiSG8p8MTz54EEnjMhS499U3O4Y25frggf
9OeVMW5ss4eyfmlc0Fw08HQqJnErnA3nyeK8vrqgyI8807/Tex3o/EqhtYjD1A3O
/0P2s8ZowqrXgD37LigDcvzUNBcFIEJIBilvtRPL/JLeWQ+SLzYQg696DVqWU6R1
2yKvRjhZlq/yN4ThuPBJcngwcu1LFsOf5BbPasoMsXiaOC8XMPVqzx1uQ9q+Ooz8
MIhwDxuRnTEbn39jlPxsXD21bY7PCBG5lAhhBqI66L26nz0X+JcBJefDmFpq9mki
uev6LoPXA58m/IKm8x4RNLwEK6nN71UcfYsmLDmgPD6TiOIMvySY28BTygPCZJ+A
tANBPxCIAdg5k3g2QS2S+2JKeurrzPJTsFBYpjwNjBPAWWSi2scpP9oMAeBl9K/N
klRbH0xD9sjrtlj11RX08NZ6zUjd69FKNJoLtOMIDuD5bhBY1sQT5TXpAJQHN1rF
+ErE1aJNmZD+2Ihllbi8ok6QE9ofvMVsgHjqG6XqCIrBrgAkw8CorH6zvba8sAR8
LeITY7zqkjsE5gvNw/TmFzYB6RMpFfTbM5gSKvrzRV+nhoN9kdWrmGFePpIACHsq
vrYOD2ymXza8dkJZY65UHu6Gd+92zcddTsGzj7ocTUrjQaRWx5fU3G+dbv0B32nL
R7kqUMOkWf6I0PFMAovTU8ekacEAnAswnz6xF8ej9Kbu2K//l3Nd5OjDe6B06iG9
yhqnj0XN3gIDVvlrkE9+Io2pVwesY702kYZh8viBTbbontQi7oB/9slj3Ao15Y42
KHDlJiyRlzSRY6fGyqXaszWHtVEZwGv7biYzkMfJMfibzCLK4PaMM8qWIO3OGoRq
+F8zfFGXeTSThNCSDBknMgruyo7da+HtZV5W1oZ6fS5xFG+dzovlDrpDvb/qV06X
f/cGAZQZnHx7C9ZDwc+6tpF1HJOQzh4Nm3ToigEa6J3CPbzwYSW1wdOcQzd4tIma
HBr9Qd8p3U6bEI2yFYHGT3YDfovb7YgJnlE9G2WdX8F1Kz1ixfE0zWwUAS+1ekvS
Xsrh6c+vepvzQtWYNfaFTHfjFY9+N+Xva/XKaD/iFL0NzqfWujxkbZD+tBSHQA2z
alJwwf0FeYO2bpaodW9sG/XBnIV/wHyueZpQgZyH96Ao1tzX43/unJIVmXPu+TBn
Ye0sTzH7txuNDlmcRWL5fRBKd/GWf/bvQFGBinjb9LDASbSlA9/NbSaPd2V3sVeP
K0WzZA+mEVgINb27IFvGsQifu0MHipiv1zCFfHOm36+Uy7yzQ+cvE6B73dl5aQhq
87zmG63SgY1RiaoxXVcl76L2Rb5CfKVh6ttAxtX9WAuR/o8Pg5n8g05ECJP1Abjy
/x0ycG/yLneB3BYJku0wQlrh0LTe63jriqcUI3Z6xy+5VgaoheFr6koLmZ8JwZLO
6relqWHd5yLiN5Qmim4CcvHeE8YBdjHF0MFqFP2RY7km0CX4xzOGpeY1JwX3noR0
UnQ/6lnY4D4/DqwI+a/Nzqb7R2K7HzRtUoGiHBZKc2M2NeKNJ7qUSQ8PESRfvFhT
87wfsH1FNXcx2DWXACrfAVsXur9Ee7tqKbigjmV4XOzMlNzVbaIw2OcGCy/wz8J+
wLK4xj+smdfRR8pcLWJwG4AI+Z20atO4ffz/1gpkph+Wv6gPZF2pNxOBZeJRSBSW
rliEe25DeqhdaZ/uNH2Zi1tVYOrRYTy65uEHcysJHLVLodKk7AyzjXe+GPrTBtKW
KNuWyaIZXB4kOkgYOzawENj5XwD6Dlf8UaIbPeDBdPtSmpH3s23BEI4VSexUjxpk
r5IyiFOge0ziFGn69EYvknjRD6MHWzCs9PFfKABTqCpymJSkWyoRCh5QiwLcMC1N
JciDH/0gvQ6wO7TmgbuRV4cFG43XDur8mhKfuLCS6gvVeooKuK7oOpQprvwIrDzE
phqiiHFrSbDC6SoUcEv4Mz1OsMRjvJLaUDDhz1QEjx4qG0H17s290XFNfsv2BZ0X
xAcYXgV+9jwNSenGtuxe0aV+xpH3ZyfWT815/3D+PipMlFI4lwtHCc62mNQsr+XK
JCkU03R+lUjVZX5nL1iNXD2v2dnNktPPZucf6x4/Anjz/g301JYsdd7EEF66I0aR
2Yxt/YaI+FXNqVBgcNLDyh8umx6wMJ4AoCci2gT97r6PeOLRFyGjH9npHrKMVA9V
p3wgOCP2I6emnyvPdkh4MT0GssGIYeuPAFzrX/sJdgIieW9u6cB3WLyz1SmT/9+g
+yQFGama0sXHfR6TxCgYrLSwRDvcKHiB0PAYcwPOFzeeoFI6qYr88NreMEWVQj2Y
H76Pk8no9SxIe2EQg3ENdLtBKm9tJOZJs6xJ7of+ibx/DwIB6AzZzKfXTiqoBF4X
tiOMs/OpKWxJFYSdWyzJqOzLZLIf85/Nlrg8kp64bg2ubd40me15kxcd1tG/pl3A
1aILFsjLNiKmjYxonDTGExykFV/42rR3w5fKIPR+2ieOuvea+IkuXnT1ZfNyPC5R
GOjCFUi0OJiwuGv6nfk3UI8I7X+U0CQjI7zYOamYh0lGCS2r70MUwpjJ6nQFmbbZ
V8MLusGdEtMGveCgZrJ9VCLJV4YjHXb/7ZEOpRhq8FGpwrFC5F+E0BTZDHioaWSB
dS698amayIX0WHz1TWeTA6G7ztLYF9d88RamhAu61sZYwbQQVGbJVv2guVSM0jDR
5ivjG+4DcZ+F5Uscgtvh8ivpT7Tz74cZt24RANws1lnJvM9WMMQWjItCnvp3t5fR
hOQsRTwr+dsT7uuw1+i9x9gzHhozdEgK1OfNd4f/fPaDxxTXPJKRcMvzz3INi4ua
kD5s/gFJG1cH9m3flyX4LQKZKZRv7LehLjOwDuLj+olO2YRA8sVOwJuu2UE7wDh4
FNES5KSDQ6ao3GEYu8taIxDUxCUUdl5GHPZGOGeqSKhgTWWfZ4Y4QQ0vvmMXKSja
rabCu2hWEIVLpKNcIB847ouxSMe0mXHFRSUhZJYsb8jgtI6KQxNYYxwO5Y1wcTvW
nXJAvQVZqTPeMqMUJdGM4J6WisXP37wc448v3ZXy0KMKNcFgIU+CUGuLco1CcY/m
g9QcsMnD0YIjqjIge8Hnz6H6vqtEMgmOFOIvl1sGSUPeXNyZsvyxDP1/gZ98Cmkm
banMYgo4bXITY4td+hzjyUgn8D5EggcAwqzqAXhGurQoIEfDMIZ55C5AEj3CqCnB
ho4Odx/Fv82GVZTGMhfTGY4NMqVmLy5tuwJ2WbVmIryD+HfHV8PbBAsA6WQ3cW4X
m/wmTanMVPrHtyYIlcibgh3heqneHqPuVnlqYPKTu3TFZBYmpJWFw+2UK463qTGp
AikBMUh1l/8UrW3mr5ehFUnB6d02JS4dql+nOoEgdjjBsmoOFCbLAjod9fnBXc4n
flW5veMHpDBIpd1yKezQv/EZ/iEBA10SH6n89Q2Y1YxH9Qf+96bAIL6SjMkIYAMZ
AUL5pNmaR18tB3OHfynqYTw1TmjC4jkXzTMBxnBQPduiUfOtGpX6zaQF8FKCboCy
UWixduTEifaONGlaXADlpLdcxVMSHbiFvoI2IK8+PBJsRo+NOCPFe9275KKT/KdJ
rUnFcTDTHFtTYxQF0zOLsXpu39V14M1Ky602HxX84Qy0/PFi9sTL99E/8GjpnTxR
vSXN8ziSaG7NBu+LNPKukRgWaEnKDoy86EqqFmYMsFf0tTsjZPeq3yUyMFnpMzUD
/VF3HCobyY4rpKU0Sh9i+vXuvR3fYK46mH4euZO9m/uYUXDYmGkFKeKJmshlcdd2
qqWbF/ZUEeoAioFlqWC5HZTgMseF1zZp/jN5EoGEOUCVGuUv3LQVu3fcVUJspD1L
wicmikcPdu9j6HvrCp22DNasGzOiVmCaYopPyxBdUKZQbzMK00qos7Sr9jQgCzEB
qHi57AXU6Y8Z3RNNqpgTFtPwpM7zQvmFVkSxF1I1Sa94Siq/EwnCBRD8H7G4mzje
E2crHT8mO4x/dofRmFIIbIrLWbnu65fe/2MDi4gc6j2zf0Yxf/bVqrzzVHcnqxqJ
j8Q8WEaxd4Na1ocp5yjFOo1sk1iC8sYfF9cPoLcjXJnSF15Id+NQltMIQ4xQkv0u
wiKMw5vDxNrN7C0ZAzb+y4rpIehcb56IFURAgGSIUMCOT/7nDJlm8Auu9wJJuNrQ
d2gRMmH4VhAtiHqbMr+g71rtvMWyVqJeqbE1rBgApTo6u3kevM+4TzLNc+LJcqId
uczboPPluq6wKASgXu0Sts0Zzr4SctksXAaGnM9iD4PxEYymHIIMaStaQq+Dgk2K
skkw7exy4AzH8jkFfPIOKLB6RopIjMBsNvxreMFbMz5q761+RlOcYyt90rG1QTto
XBaKMjPKdPdPGH1vSeF5EdB0ObuJw53jpLwmrjfy8O1yVFEms6nh+sqTYTCkNkz/
I7TxTqken5XhlqYEx0mpXWBUr0xPHVz0Lv8c0cQx2tU1BstM5m/2sTxqbk1OSf/j
4eYvwVQ83zDVj1auJTX4iXkKPst72oGQelO3tna3C1l9FbiAE0Z1BawBrCR4KYT6
e9lam82X4Ol7rvahptBoJEF/W7nOrAslbhmWxZE8Kn8HXjkPxMt7k0lkyWyk8cel
cHjYh7tH4+ebQ35gbG4ZqloeMSbk7ycckVM17rTQbznTaKgWe7QxzHGTO8PvQvmL
AK9QnZ/o7CPbg204kGD3NzdNIF2U7ItMZwYK1EqpMN3+vAu4Q7zI+UtywH8LDpYv
eZFsfrreGS2giT1q+TyHdlIYwzcyrY+mBCCKPitsSitJAclUclNvjmqGEKo2KaC1
lYfI7gYwXq/jNBf1tmfZezvY4Uax66nWocwAJX0H5RlNbQ0h4UbIp+ykyevPNa+N
M+Ojq7kyNoWJc4YoqIHhMn9XXqpScCR3W+crJGTlvwfw/AlR8jR38PDEKukB0+TL
gw+oPgt/kce2OzVZdPla3ZlZ7rkzGFYcpx2xikbxXGc624CwhRfVwp+iltIAHqAE
fdZsywKqnFqshBeh36quMK7oadQ39fd42M2IEG+Q8RMAARMwNqtxEuSHqpn6neZs
s5uFsY6i2Ky0KHeip9P+6Aj49YPphwm/JaT1uR0sJ+64pMnR/d708uCkGdrG/nQ8
C4PcAESnCbAeGf2Zjbc1enIj2uVSRNiNvfZ/fGiM/1lCoesN07UL7R/rM6C+mb9P
8p51wYrsnKYf+hJ5TMkxcnpjdN0h3YrPfaQP6MUkrVkXd2JzgEtAwRwg9Ba76DLm
H6EF295M28lDvHMiyu+fd0kgPM7CFQ2nt/bz0LKtsAQ4D3nDh8IFhgSs2Gb2+1wR
PfpAYs6/K/xKPs9PZL6vXn4yM77nAjv0P9WRakRR3NzrOKNQyxtUfFXhOs6ilTPh
sYyvX5AsIrWHX88UKPGUd+jVXu82ctJO1yPtQ8b7MyaKB587htJl72MFEuul0Z5K
sL7889TWNkEFMqmVvSNyRrvztCNoOUUjKkAh+ajfoMAN95IY97/Qebor0FSYm2Mx
zrHGsKB0ucd6OJx3rw7Dym2avs5Kppxm7canFrtBEDNfKTxOGepd93Pfp5Rlqf1a
NX1dcK4/BVvT8KcfLdpXfs8l2dSBw6I3ltEslCHyPE7Nbc8E20g/7LEwUVUtp4wd
UoBu+dmVWBEwTmldmPYg9Chlmck1WMnIXEXDRIWInpGVPX9nOg8n5rblWCDmVFJZ
L1R/+MtFtGr1HuuajUkA2AhB8MVQQihwFhfXrw6ktXxRHcT/uieUn0nEp4MmEErh
IIYqJCh7/6U/1lmTUqQEIZJo0CAPUrpSZ7t7uax1THmgQl97Jyeux3i57601Sl8y
ts09l50HBGcglGE1mJCTB12CKaUyth0tC1NLxFkCVzrOX6UmpTImdTKyX1hBbo23
Dpvdm69+lUFxWNda5MtXtlCa0tJeYj1mGu/OOY0VUpAycmDtkCO3r0Ut83Rmp1Vr
9m2BU+jX4rfVMY8vc67QNCriZuayUKzWixui6+lTA/+1AjgbcsRsdqDim7+ZUsNK
Rva+MXDRk4Y96T6DlBWGpnijOT4MS6w3lTLiLGxahQSRx9nPGgpbHGpT+2s9a69x
bNiK0VKuASIKpN8gHFxs1f/pAh8ewLhMQCef4Jcjevl9oXq/k9cfbW6zNNnwibXp
y+aaY2x6IXU6e0zvuXedzwBowR25ff5P4gxglluOpIQOt5phC6XisiBr/fcLsapv
C7SQCuk/weg2zm98C3PCr9/rx1dhEmzj6/HoNt1snLXv5veDt3zRRyDC+twkCeTj
z3wDWjPEIxarfX1t4eL3vf6fM9xZRP2X5pcFmK6UjWq5C7w/I6JGPpxmF3bfryzn
wniwwl/1TjERDfK5ikFno9rUuz7L+dmUn62MNCQJTBBRnwLXyoPrsN1CXacTIMzl
74Y+ulhU3L5lOvZlvAuCTwoAM+kNBuw9V9K7HUQH5wNsbKm3gFJ/0JJ741lcsDBG
VYIpDFrgYijrF4BYHxX5Fi4SCmT9TFbVfvHucSwStyBHIirifGeXUq25ZmVf5J84
G1QcsBhWc1CNzKfsqDbBqhBMXqayQQSGrEMy9UxrRGYONSYpcXrUQG2gcmGBAgDH
EdudqadstspXpMhCzNvICrkWKoCAvpX/jjzZLfDPrDJoROCimoOJ0S3eqcFMDvHm
IeYv4njsFcwRmN6XPTKGuVKHBURiLfo88oXn9364c9AQy0pngoUIRcmy6ttak0MH
/B2EWOAkszS7Ar0QL70IYpiHRINDjHcFZfPXSinAAnlxWdZtVvnaXCnTjFypiQZr
q05/kRWG+UDRA7iH9hDvWVzVcR3Oo6vOWFa6X/T4aNfxSc/4P96Wdgq8fP2Gwg6X
v4LDKGVPEm6tyItodhfFzCdwE7g98PvydOWpnbXIMeN8RWV9dZozi/thRIIrmNFJ
paM5ReSlBgmZ0Zvyu9rgaqGrzKaQm4lxxI9xGq0NkgYX+JBghpP+mjlcmGZs77D+
TGW5BH9oGVsj40hRUCGRWp/Jjn20NdEHp7VvafUDql2e7q23765YDsZDO53YVS1q
YD0DtNJI0I1Wz2+w9NIkPIlZPNvncqzFlAjvHC3LmolSDFwKB0Zp3Cr7UL0ZY5oB
U0JiAGWsh8Ue+4kUIfYmnSJY6jxOuhQ7GT+hxdy3hatwRVFoqE0927eGvlegl+Pp
lXZp30bqmaZ6f8Q303W8wbUmfdSb+ovpagNSlSl616u4SgLoC4xuqZIlEeVBkiVT
tU6ESH4R6tYMXPa90Lcuc3TaF5byuKR3I4IES1YFjxjicduaR/GCCU5o7kgTP75r
zzq7hp6Dub5WitJ+iMzhX/Bj+SsYmhC2Lbqsg6f+P4f/yao/jrCqwvfFWOpWshrG
Tgq3aSLJJ0Cybyy1q0fecrStUYmat6JYdGFyA2kE8H5ofdflXSvG3s/AKwp3i9/x
+t4Ln0kdtUIXFt8UAkfwI2LwUQkWAKGrTyy+7ZyviOkQb0/+8p/fmKZwFLPx6t6a
SEIXi3QjvONKtHOPokbFGrUZ0D9DA+tu4y96Qtjnnvakzqzk3tVaQEaZctzj3jf4
MuhUi3SlQH7WnaVndYApetYfHZLuYYyjB4x3t/6gtpvxT/9mxydgnvHF2eX4xY+M
s+hV11cRPNLoXkpFw/lUkqnuFvay2iuNFrAQZDlAS7GE4yL56cU3JCWJvLmCviiW
t8Yn9IdvmO5ClGZgQ6AMtIruQvPq8r1ylFRTblOfXrXVmLWV9euIYmLZj/atsXcM
4khiPIAll9tY7ejLheFcEdim3gZDkR0RebgWnO8rDMc2dTxXK0R/Aw7MJn13QPUx
Io1h7sRPb8Q+uQ8H1iMP90zU3MOFlv6cFtdCHyYwrr9DDxPZHnEZhOXAk47JMQTQ
dagJ0pObXyZ+xBgkJ9g5Oh2HFIxEUicoHwTqrRvidZ+DH4OE/HXDHqyzAuLcpH/A
ggna2FgV4zOxyrLUEPz9tXrT5+9pexP7u1PSyccfQvWxo2m2O/WNg1WTuKi0Mo2j
A1l/jaziPPTjbFjkPeyeIfQyJ7pLga82jyYMt2uttRrpI1LrrXW0sBUeWhqv9kwW
HkBFkRLDvpaiFYiUMX//KbJ2qjpDFWITicUZsICYSLuYWzWo1l40O8GDj4RxUl/M
nfjCMrX8ohjR6ZSq6dNn59kttPHK7DYHrTvNWACFsEkkyaBWEyC8BQ49m76xbO69
CU3OXqeALbQ0VOREF5EPAIQdGnTcw2DZ6IocMw3wdmWicGCUCz1TAhDmk5g/eVR5
enil305eb/PGKFp5Sh4Ae0sTss8GTApWdXkkxpsj649DTq7wRRQClyMPXBLkglKg
68VbQAj9hN5dobJzrEeKd5fyK87Y/kEGY2TZ+X02mjHdQOg2fLXGo44nxtLM0UCZ
gdEWE8fcY1CM1SWxMOyuCguAeZSByaSnSNEmcA7LofqWa+/TjGwwBPbAXwGrFknx
KAZf4qMuQU1sjhmp20VJVOco+ozifBw/Aby2G9Y8rA4XuofQwyxDQLKsVixGZJU3
m9I24foCqe0uOFhXs2KjnPzcVbTU8h+PEUGLXrv2HDuZ/Gyz3fTSjr0UJt194Bxz
yd/AzM9nmf+PUTchkuaopIsddsp3BhHn5us/WLFxBt63YAiRynlDo2vM9A6kSQ90
YFz9EpWR3GIV5mhHkMZTYujWRYV7zb8ZxcHrlG9dQTBJdE6HkIVQvtDcdvdJ/ZMS
WZJomAV9jep4jZIuWkPLQK0gGG7yZLXgDBB0A1T2QsX0XrFUkVo/LjksCa9RrjSs
jUC2pHHMdDnoihNbGrzw+qZqsFWWrAwaY1u970l/7vkt7LOWSj5paSSEG1L50Lys
tWI05rtYfsLXqGwvnJa6OqJPAGdkPNtZLIyAfUwkNY7Q28N+CPrSCODiogh2XvEs
II0Xq9cquO3SpNCoTselFmfXF/OxnUeFcRYGMYiLXU9iuNAJJRBq3RopKi1dk5DO
418G2CaXA4VGl0enu4KzPpICi+oo9iDeMxOrwRhKGqv2Y3g1GN1W8F2lBqwu3tmr
jczKBw7Zl/fUP7vmScX6khWs81amWNqHYkYdWwTsKQKGYnAxHJzxFvMFaeKq6Ha+
CxCUlSrtn8iJ7f7SZuq6YnN+0Squr4ryVkFPMP/DdYcO4806cFEQB++3kj25DtCM
yXHwwQUF6DXTjB27RyI1Bbp+c+HLHAFbrCArff0oWpCk2mxOXnmiV5DJtebkJwJF
C3aaLKdh/FIL6fkUiitiXkaAJhA059Ve5eqn7Q7mz3AMz5d5oeahOOx73Nl6mT24
3OBRPhK427d4Fs6moevrrVVElLDCUjKQ3xsz5VBBfOIdsB/AUzRrUCtubg0mQHp+
w7fqWC6hJsSrQdSm6iKugnxJNLYdfR4Bn+Gsi/BsWDbDEQfREFOJ2aIbNLXLQuc7
WgZ3V3TWf08EzNJwlEzKzt15nnMEGZ/mnpyLdM5tXTPe7ry0Bb4JOwaU4hwjcYK3
XQIiRwc7q/YOEbmpCeMYo2CmFjOl7wohMP0E8IpcDnq9r3ZAu+eJOlwimKUiyJhL
8lmEYjCkMsf0xleqW1M3cBTG+QPppGJTwk/tsY9L0N//eDLcg466meUKpfy0Gwj9
Wg29VRi54qH0WuwRwxxki/JFfTpY3YBczeYEhcQ8vYw6dZXAjTkYldk8HkkkoUQF
DBiRuzDkJ74lQ0D+UimI1nE2sDVNOVo+Ydl9vAIVoVVr6PFCPx/nmbFF9Q1K2nsV
1ZyjkS8I0s/Cimu0LiJQy+bBlBI2trLqG8AK2Z/yEm3aXekrR7Fjn//9Vyb3wxYv
9jg8AsXpPWxOFNeYAftJ2N+hqq6iuaZTWZ10mlLiMqHT93CeCq3SzhonZq3Rm+KI
6cBfaO8HLoBV29jrVMgx601Ee2WxrR+k4zHGBLKZ4bJIeqSDd1jV9hs/4e13qrwX
ydY1KSanmOh2KLF/UQLSRtLiwN4sGp7fX/b6XnRnwTRv5ntGngCJdw5vdfGPeoLM
mZnYAaKPGTARZLEj+r7VE3ZfF5X/jeWrCftHWAv4w0cWEDlUHkFTaygdHklaKTI8
i6xhQWZQwc2b6RMDVbYeFiFlmZsPfXTsgQ8qfSooCbLx7D0ZfX/EtxIsD3V7IK1N
SRdx4SzRoneTNM/svZrGGImjl/qVCstX1N5kjcSDI5sftYbiUMgN81Q0Aslp88wh
AzlxrKzIzW1LH5IofScSJ7co3Auvr3X7t8BSj9+PHlmr+I0epqbfa3OPAfjCBbR1
hstrrqdrJveZYE1QIOldSAHMp0yAfSW/BqONcxdHaAUl8K8ILTCC8lY7Qr9U6rm6
fIJtLSn471JHgJEha0Kh2cGAD/I82VVpV3+zUhvUqq/W/4B47jg6xyuU9BeyO/+l
rQZhrGfsneldtW3pBWSrCQOwT43WppT4ExqXAABx0Np4GXEBl7aYdt3bvMVO/EC8
kfVGSoCFFmW688g3DYhm7BAHYBXbh4kc5XQZbTG+YIXEYH7ZAZkDO/FhjzOfrebQ
CBITHWp4eFhy3zoErsdS7iFPTubemVh9Cd1Og3lqDcrmpkIbuoMk+fz3EkgwzgXZ
8NhYiX7iVesv5tQylviGpMhqwSP419kTqa9g1sQ2nDdhLZ8QOl4xonoHm9O61Nrm
lG30z6QO7YpSVV0X3j8AWs2g0f/zoPtni1pJFqOOgCDIFPrOPqOUytqDV+st/eKz
ERDdFWjXX7MX+v4/Sr4l7n/KpnVIsCigk/rz3bwYiaFmMFaWIy2Y7cKF0eogm7OY
r7PEBFWa8jwI/ltbRN3eSIXVu5G0XDQGmTg1JuHQfrPKEF/CR8utojZZKoHER+QM
vn7Z47agi5sVUWT4o17H54vkuE676tBPZOgPb5mRqr/UhjTjmiYSMbxmk6JI+Ns7
NzmdkqtZj3JSCtgv8DxsNDsFn4lJfkTN1cjQ9BcVlJJBuybKuFiklxGGot4NDvVS
EAzLU06RNRo+iiCgtBa8jcNOlgIglzRvm9uuPZVZkiTN1AAqpuS2E7YseSR9S+Ue
6++7rQ5N01XpX/O2lTj/P8or4aoi2MsS60pq6nvIrKCHS4E0ZZHptGWS6u4e87IW
vzqKW9A2AhOYOGmXalLnC89tR/DA1s+qT6AjXE0S8thOScFbk2aTLgsyG3MqCy22
qK1zSxM4BdAUIpO/8QppeoYwLITQfwyJ5G52XnZPgstCmMW5itsDA7FuR1BXpOrl
GrOrpX/RcF9M6ABgShU53GDfVaztsdpKNiLrYBIgrHBfcy6c0Lq/puv9YtjSihXE
3CXD/Y/51ZLk88P6yOVlDahaeC0MTr2hOeKJ7918RS96VewT7w4CdxuIzJ/Nsri9
CO4Q2JvPqF9ugIvZfnRtS7j1FYvvXhpBquFT/cO09FjPte538Dx/ETL95WDidKIb
dWWw+dfsutFWHUzktDnry9osrRodk1k9u0Rw4yn6Ay6CNctuE1pmAnPZhj8+sUMM
+MdN0JcqaC7bvum5LxOxSOtcY8xmvdqYcpVEV4Rk4RAadW/YE4ZOAe5kjUY15/AJ
WUvtt9NppXgIlB52nfP2MsN/d1vZTGEvOCaUs8MaYxaWfwZsnT1dQ2xvzcyZxmVW
73QRWlxGIJTM5m2L/lwjvwf7V5Tp90JN/jiSiddWNS+BHd1w+2Y8TA8R5O1qyxmZ
2l5S0VWNi9kz+8OwI7MaTEW3F0O+7IIe5aFTwcBFrEpCCfbS0FFEpWGwKkKZZOgh
WVJRr6iokzsT0VxP/mytUB3b97739K2KUN6J4GBVIKgQWnE2f4+23PCLJQmFYSCt
oCzuMlnnz9hbJPscjkyFjpajQArfcDHRFzyiiv4IYfJjpS34Znif6XsQroNkOaQc
fJxXZtqaguHw0dwvclyFYpTm3dhhdchR0Szej3LjjPNkeEyAyTowlHuy0TrenLYd
WlVR0Pk6RqYZApXYFM3upvwqz4wdxEt68ydPVW7qIAbjRrW6EZs4lUTZelE4utad
3ybg7njBuqnMOgpVA6ZDUD5y/EENTpJiUQLBUCKI3ZOQQ8L3oUutlVCyuMkbAMZz
9Jkq+YiS6AYWFnMRMxZUSeL3w1mrzVLfhE98JbFg8QW6cfjNtQalS2NIX2xvYvjJ
uCuDSK7ByVIsRxVO1iWOeFQcfA0alonlfLBQ+cIOawZZR+erTPcJpSW07W6so6y6
eZbpzIcjE4a3PrlooaY0qOky7W3QYmtDYoy3JYDPAtKydFmfIAooUf9F2G3YPix3
Nby2jP7spbEXg9FrJlenwTswCC/81X63LsrjYNCKVngJDNgcxEegB66M3/sWycer
pbvWAJPzVcPhAcbCFM6Ihcw/+rL+rDLWB+xVZlFpv64Xj1npOgo+fDQ5VBQrk8xE
f4MK+QdLJlCh/XkT2jKHciBzYfSZTYK/QgsN67eg77M6SgdaS8kg3MLV+rLX6LQ3
gNZXoxggTe5OyA8R0KmgsgOieQju0bao0Xli8f9zyD4NUtc2o8MgEGtJ8PRs+lR4
feg0nUVXayAsf/Rxm28ujN2jAvQLRbA3EwG9XXphDXLqnbe3k0vpdd7aLvEae8FD
UEbKfwc1p8g67wBLeYt2EP2YYTIEsgCVsd5C/iG2ZZbmPjU0eGRv8gyeFEvY3Il3
U7FlSlLJRgKBsvBZfxNS/50OJe8yVaodidwpPb3ymiVR5JoK9DE6vz4HjWAyLVpk
UGlKxjq4lRr5ZeVPziZJcfASmLTykgTMvm6Yta1SvO3Tx7PKwK725ljliNXrdhV4
GV5H++vUeV+W3WxK1vHKEf5xTUuzGjjbojToxlqMLW+RQsxR/FOwDD+HxrhYAYMY
YPw1Ukb76YOQBAQDln4OzySzSWvanE2EPDrCtUqM7kGmr+ayAgShiMu8XNPFX0s5
4GMuTxXb+qn87rR1sqpU5C312higIU3amX4hvuvUolNsJ2u/RXWBy75zYt59Qkx3
lhxISg8K+HwnnAmEwkrK4a60ltPj63L1sZT+sh8U//CXyqbCT23CTDkBlY2sm83t
kmvPX8q58RsJnYnpKZV6MPpM9MbQ3Dnc0Pp+1img4KUCATJD105HBQO9dbPEOOk5
tzsVwbHequApiIRu6a44YsTja6P4yTMEZzlZofBaNCvz1Kt+C/IqhSBPXEdv38Oq
CsRNBUAN54X1ULza1d+C4a0ehEQ3HbdX44qYHh97dZLuYOn26UKh/PA/LM+npvRK
n+Rl8j+1ixFw1BYkWQFG+bix1qc7GdF+Q1ZtZv5hSYVc/Zo0frRXdKYiE5Osz9Sh
DC8NSlUFMu3XTV4E1SnLmd7lI83HH01jy/NyHjTRw29GKcJ2HtGmJutsFthNzi7P
TAjc/5ieYp/I86ZNSUtej7TGgprFjhGDS1AbhLKT/2Uw2+Zyd3s3465yvor7PiTt
g45vTG5mkNGpRfB7rmO+qsQd704bBxV2az86MYmW7CdjV1Q43z9wO8jE1KDj7Bya
+FX/0b6H54FxWcIwjKYWb4T/17w4EjLnfTA3sIGrUEH18Kb3Cz/CKt8i7mST5GFL
Nlg6kh6Bl91fNEsxvr+FGKVs9FvgdJIUZc5d/sf57MytsQz1dAD2ndkCJEXmVqB3
lfk0o0hOzQrHfdj0g5AuI/nJZNGh4vyKaKikK96b+v0hGa61Wdqi85sVlb+i1Xr+
DAkUyDB20zadbsFT0RbxmZ2XrCrQb5KEjmygmZYJpE7URaMmxVFggY3+zSL7+1sB
WhxLeJfe+TkGtnobqFQRLppHBroytYS17LoiPNzipfvIslF/pPd0apKB8H4H7S4t
ZsafCDTm2VprygIozuUeRCKrtaAnmIw+tQvoKZvCsTvnc6ke0BeSwx994jJqseDS
yUg15GEGpBoniUJCjrLVBk3Hr+wBT99c4+lqm1mIBqzhjx1vHjCcww8jmkCgsPxa
iT8NHCshlX6KJP3pYDk4TPeUUwUpogDj1OJJd9YFD4skUjQo9qlDJMw25TG7fvJD
FrBOnAjhSUMJcYsJkdlp7CtWDbXNRUNAC1vkpeQfbYXiizmFWOWClpZKpvuZVqez
VeX4EXXS7ESO5HiV71IOGs9ZitmxwSG6yCD9oDnqXxZvomr0001IhbRylyr8JsZ+
aNjTAggx5jtIBiNqzJGqTOCtNsczmS8GUHLppYEHHDPJLSf1Abuhezdkis/xJdHd
ir/NUov7OfSSsCRB8YmX3k6bTf2uaJIjBmHLoWS+NEvfTyxH5qPW6nrzo/nZnEBr
wppd10cqniJ0kzhlIZ+U7W9OqO40qNO4dhpybD0zV8tNSlZANcM5ucC+AQngmEwQ
TJNHDM0cLJA+5TFx/W8A7L9Wi4uwT+6kCxkU5AqPPqd1a/v2nHEz07stRfbrOafL
40zJwtypMTAARiJMnNg84+9zFZTbD/4eaOimFdoC0eujjqxRatk5c3bdMaN1RVUW
zmm5yNXiGVTOLCxteqy2IkqdI7q0/eOtKd0fpItYw1PUeioNXvpxjmFnug+Di48B
xBJtv2oJRJ2Y306lXcI5EQvsMxIgkZnknPUVGtzKxu0Pkb6mZl7v9AouVWBeOLfD
zrMELtDo0BhEpSaffPE+ZkhQ1dw1qCT8DgXqaJeO0eF6V5ajyi+VNv8vu6pVQtte
VIyjtt7zTJq70Jk6F6C9/zyRwH/AbURB2FyxqK9ZNc321cTfekgMCIXGY5T4DzP+
5PWmNWjYMv9HhLx1oaQPcx7vA7zE1YteY6goF/82xpV3eRTxzFSrIh/jreuUlYyg
WyA4cqczWoZMEgYGCtVNDboknbREeOrQpKbyl5zDYGD4vGFsl0re3XCW8L0l6Y+c
T+8jgwkfdMzUe09JHXCEcH522JUSk9VlgZxfaSelso6XAo3XkblwWKj+LM+kd2bM
+SXlLi5d4IggBgVvxFHi/OMOipa2FfYgGnOyaQO8vqWWosUSXP15ycFs28iY7z2/
RW6BVad7oGVE2oLjj6Xia4cyo0qjRAmai9xBvPfU4MX14yBCKrAecjM430xagTVT
dNLdoZ7VgJZsXnUtTeileyb02HSFKCSuKXNsbbz2Ij1WmcqDtV7pRhCCOavDqmSy
+oqJSdec3MAD4ZJ/F10IE50ZSiJauBi4WfkKFT7RJrI5MUcvdHh3ErDWBbP8e4wg
RMXlS7KHgFoKpSF8dFNdGEpzAjAaYLtbize2fsV1QdlP0LKJ3vjMH5zd2vbAeOnN
mEjxgGWhHy/dSprQYxPk+szbBpjC8R56RuNSdEvKHDtjG/ey9C5cC+jvn0/oOyKX
IVQXuIqYR1ZrG6CkvFbrVfzRTRGqC+Pwam/2T62KQiDLxzNKLYo2rW9v/abJlyBG
2zKW/lejHvmvQNcT6LznvqI63QNyXA2o/42pbwIUi/k9mJPhEhZvrvjeWacrMhY4
FFiTmcaFTKJ4tolc2R4vd6ZefNhjQZMVDQVBISe58DfC6HWFXquEZFg2Zu1wS2Bh
qTimrjOHdEpS4KdOiLx+xBUXox37NMqwjKrDjYwCjEfpO9s5DHt8HH3Krf8nBvU5
HtheCbG5w5N5QMQRqxtcHFtyKCtWHwaR2yvqSL6T34bNCT0VmDuHj1TXJdrfKwf/
rh4rQAIl+/1HczMjoyM1cPY8ow9XOuThkA0po2FvPUSarpyX3Qt/M/JlWKGZXovO
knYTtTv4wwbYKFN8tH8lSHvwrHTuLCUETfWYNfbdtGn0akLs7QFqWjRTbAUn20pX
QNz+pmKlmZox5i7FOxgdu/cYw1qEt5FD0yOzTEi7hhbLgWFHjK5APzK2TFem3Dlf
GRImNWTWHSTLpVEWl5fyL6kfy7HCU5SHQk0QnzokH6EO6inm80GR0W48QdOPq830
YwIqJmpsGdFRpH3ocjHZ4Xf8TS+gY4G9JyteF9RcrFoIyF6M04bvtymaLH4e8iFF
eOe1nEpmLW7gdhEvn1w36ECc+xNWtfPzAaI9C9jRwF1/wSXOp3kJXTwe+ZKlpVs3
tnemsgFQGMV8IJclPc+91umXw32gyzDYa0CW4laLJcQFDiZQPALl/+inpz1L3lqC
gTUskmgo6q0O7lBVgNfgBTo+UPg8o7OnButEy9LhNCU0k5UFC2MVB8HCb7ESAkU7
GIomLqK2Fuz84DpDCDw67a6EvMyXD83Yv+LaKiuxD8gV4lUwNnX2dweFGl0dq5c3
WMGb+JeI54J/pAH1HhUc12PVLddGu8obxPnIv7HPBFqmnXvMZhBpBjPb2nLNnttF
a8nMiYqxk9xkjzoD39zWwPrmy34iEPDQXnSFKocMAuvaSIzC4E3gzQu5yUClnMLi
Ri/l5d+GfmOmv3qYFJOK5BJrb/50wNw2ywxTvAlnA+fReNTxmE8vfJHJ0+aearGC
5HWlB6o3q2acZ87LdvX/9qY2yAwkAJrL3vc/yh+4myQIav4Vm/vHcTBd1fVpSIyR
Q32AUIYrO/cp2UJmdgvI1oxbWqkpx1q/tLFwCeQwX07JRSPf3FvZHsne99ecjdzL
0AVHB3651Bus6DRrpMuJvTSa7ru8MUgDfHW03YMdSKAtD4Osiv1zGBcG0WegYZ7u
Cw1BckKnsw+7R5A3eZ+LQLAWHC9G3YYg+JsYqDkKymwujfYxubqVj8ByORRdxzdM
CH3t4GEdB9edjS3iUMVf4cPp44sXwK3wKcci76FcZiy9yFLojceVOfD1g90WRaSQ
uKGvKMvu3mKlxW4lZhj+SrG61MhDKNipHzYsaxHB73ZIK1SU0fq1M2l+VL36NXan
S0nOWaOhE2IrcS6rdx2UfrLjQmBqWkvcuf/X5hbdv06VcbAkYHdf03AF1/DdlPEM
ERIafIJf/kedYSqC1TAUIeY5qdXRkEOYtjyvBBqUdE+ZiymH1HiiuMl8zIMNN1c9
W/vvw3vQzNsrWHjiZ9hhXcfDUT5m5QtmEMcqiqn2UA9NmAmVCXgZzpyFtuM1aE5Z
7qrJAy4FhTs8EyrzbIQGKocAIw8dwKahOtrBtfr2F7g3pNJT/kogBaiRyNngRbVv
CNlqmCrC4MdIjpH1jQn++/rNEVmnnxFxMMXjljIPaYD4w1gM0hNv2bPFw1/UdlFD
jLODJj3DebJfUfgwpeJSBcb4dajMSKFlcB+BSDBsnXA6lxWBJHB1PWJDohC4Izg2
FeHB2HGDG5gb+zTPumlUuVVnPN+LgZPxMXz8Q/pEso7VyVQNNCOEe0Q+IfOcJYF+
AfERTQmMYDW6j2e3BcZR5Y+ikxR3u3iB3Thw7kXUr34M5ELRd0MoP7wcna1kMu4h
DWgtjV/8/96MwS/irGdAIDT1BaHzITfaoRLgL1Ao/G/cHpna7n2R5V2MXl/dhISG
kPmvEkI2OOb9CueLoaUhZyTazoh0WKy3EE2n9XKRLL2T2v1T5yc15IGhUd9/AcPR
r3WYxcz0O/MYMlmdpeWlBfUneCwjDfENvWWVrJdhYs/uFuRQONlSTHlcqPoZ9lUW
EtdcASELaapzkA7DvAj7YczECyJEFsBsMkLAQdMXRb70yWi/KGVReDScNzwKU0Hv
9xfN0v7lQc9qMlJl6k/2s+bxtJoxl4+q3AdqK0ypEVUe4TheWPNoPcSmK9cI5Xjd
wcWZg5KcKGbHMa72sWE76iyOPZBkZWN5aQPdjClm11td/IFw36Oh6Bl77PoLaPur
KmxYlQEX+IBGqz++oh5EgdZmywL0iyBhPp7X7LVOMre8LQ/ZIWsA7MY4vKxXiYmN
7FV4AXj2j5rNgP2vdbN8v/94LcC8uW4rrFkU6I6I2kdu7q4oIDlqGoUgm5B0RszA
UefuY3Wqpi8tRAuQESWX9V2tpyWkWKGccbnTNBBueh6dCU0/xFwDDkGJTWei1RYU
ACcc/h7503RSot52O+BiD7Vp7BndnVjThtI4CK30Ygxb4bAqDbzO2A5Jc8RTyRKQ
AYZNhiikuJK/tZehHdj4Tg5PNhKUl3pdPvLENQbJYS1rJl5u8I0EFeiqzBrIhrcl
EFPhbTlPksdzsqXbbsygx9MpjCz3CmIGAz+ngBXwc589gWW3RH6cCwmcJZCzgJp8
18LyoZA2clgdIeFVlr5OHVvzsvsJZpP5keuRpA7vYaQ6fdw6leOF9HAM0BEvmkv8
OVTaCEkjP0BHUC2//2l6xOjrL4qhe/aX9skjMOAwJRxYUBNu2yOjsRTX4nAohn4I
lW4ZPbLSF0o7lOxozJOwzjZVpL5Y2fTbs/04fyzA2KJqe2YSdDGRQ9wK57UvhWdg
E3OSCeuKLxnJIDv8IxPP/PztQG/Bw8wBY+Zoz/KzvL8/3+8+izOYXU08mr6J66iT
E8s0iEBzLz8sttB598MLHRYGEsKS/+mRT3e4y/9iF/OT1/ZXb3GJEc4WuNVUKHgq
JTNQ9nO5GjWnljE5Ev9s2Yi46tVscWpH7SuZ+Sm5+6r5heVNddy3ri1RCES/HnXb
Xq2nl4/uzAfBH3e3LccKo1YSpzO9oCh//YRhD0Cgg8s+7X5NRXvr3mSc/BAU0yOt
yu3gafZqiPOlwkz44p7JorWvD8MjWevKXZEmUbXXf6Yple90N2IzTAO3i2VbXiJn
55R9Fv+IpBpyv3K3j0RuH4veKUpQ8RLRtrZpmV/pv6BthMMnG9dIMqGrLmkQA5gN
cyMeZgTB6K28+TtHS5awDDVraMnHcYupbKeboxMtZ+Mos4CHtR5wgvYpCGT5dU/E
RdxJVr+EKafme4g4YpDfp9/uc8nRmf1kYsvGTymY2Fp0PRpeToA0rSudQv8GIA51
dRqb4n/sIgOF4HP7px88d/yW1LGSpe6gwtABy6KEtlJ9T0VRV/9Jw2yHpxfQRhi1
nb5WV3KpuWBnIxfwpwM9Uodyv7QUYADRws1MFvMlvBT81LzUueuxMtABCWCQ97qo
0CXjaM29Qo+bdRiX6JY3qczkhPrnsemZ5NPveBe6hO9CTn+V24CSpmNWGy4QkJxT
MqtJjRV2pOGMq3GGYHzFEhUn5E/0GafpKRvqNAb5DPsKBJBoqGBw5eIKX+DmRw1n
HT0i8PtAExvglW1ePS+9NazUGOWsqyutAPppkyPat+oCzlksB/YXiRWGZ6POJ+O4
oV+q5XUYVzCYG/Sgx71i1vAHVXHDGlMAMHRVYtmxlQQj5GOcwP5a+wCs7CDGniWb
tEdI537fKWhqK6LMOY7FQ7ZYBfhbKJ8EeEKcs+Zx7NkJt75RSSEBPwoFGcHzHU3T
2ukYPqokS6QpeLNtaBSDylvFu6TZC4qwDLTTBe2pNQ3U8BPfrc40+2YqNunRN1j0
b9jn5xVPdqSS4cs7K0Vfp22hePPqQFxW940MroXjp9t+PMM3L8ssPKVCQTsr691b
IkNJXPVnWLOZkZWGI4UMxV1YzttfFPvazh/ScJyViqXZ1NNB+l9gpyAgIYHz7dVM
ZNEcvZdoalmF3ZHVDzOaZmMuVWsJN2ZubJ3gUC1rNlpxj80HcJqNvN2xsdGt8V+1
uSrD7Xc8vr02oewGkGlywfrlv8ic2vvd4pmA5lGy+QeSHQiOZJyJl+7nPVy2RdiV
pq+tYLGnWAUaN916MclXyiedI9+2fHDnqKFkTaawPMM5kHx9kpCnVMvWNI1cq1aH
H5J8/4Jw64WofPpwCrGmHDRCLLurFkG2BRn8zbQGY2UZALpy47Ow3U/EfiNqdTSF
l6+kZ/SBygG28Ppu8QGJQP2VKtKdwfGN45OiT3Wb6q18Pndk/NthbpkDaGc/TT4h
P6NJq4C9tBxNXxi1Z06WwXlI8UYZgBWZ30va87wujBiWwqNiWvlI8zmdtO21d0h1
yvdjmvFcNh/P6cHqI8GDMf94zU1T72UJB0rWRHng89kT6qroKBqvUmXM5vS0dQf/
t7JEyaa1a2vFMDyqmBnL0s5DE28U7YQrfxIyX3153muh4qFKx7zfVYUlh6tSnEfJ
EoXbWrsYescZXNtrU23Uql4doA8fZQu4Qngi9bP16uYdtqEJQD3oMiJJoOCjM3uH
sqWRZERx7uUIOh1sCvuNftTsx1HamM1e/P9wOeODGHrU6cBejliXRbDhaMAfmGgW
R5y5s8w8f9I1NGQ5Gnn3iIklmmbV93xNb15saPNNj56SeYbsqbOUZ0vKeqsBzBwZ
+8R9J42QMqW59M0DfcW6Sx6qk05dJ8eDC2LfBxzfGWnFMdBotkUWyS8W8o14/ej7
McuG+TnMwjZM9m6JoeMc+4/1vESgUduvLxNb+hvVNDX1PIkqiwpWsTfeWnxg00j9
epVnwNc8p6rqrFYeaWUyjRyRUUHuavgcr7Pm60f/BE/mqjkDIABa2UXRsS70IAa2
ON0ENas6VwFXkAx5XssL24/aE1HLmRRe5Q6wvntY7sv7/YSJ3ph7/YOwaDW+rO9f
eK09NmRB6ee5zSya9n9ICH6Ni7jL7+PnYbXP5hrix6qzHHg25hWaeNTU91aD/vYs
JKP1P6D/Ie5gzsfTYrBafexVfIYVutGOu/HE5o9LMGGzW6tI3IfcdZd9cS+atR2b
8lQRgxTPD/eZ49d6q3ApQLSGSOpNG0Rw/qDrncIEJ3dN81M4kORWjXE6oJ1sf+tq
SSCQuFYioi11OmVJI0IZpz6kQkVhgYSjhOKVHy6cIwbKdHQek9pBuyv3DUkatOjk
bLYPW9upSkkUBfmJQika5XK1XzFJ4bho/4Z0kMsIWM0NQubyR1w1kFhDfan/MeNI
J+N+FeZXysVGu/XEU+3VFnhA/nyf4rxHHHiPGa+MPb5ceXL7cnAgpK+CeaC28bHx
7W74njG6ROcMw8NjwBZ9WMVun09fsF8zre3FA7HMHMtszNCNk7FAKpWdGw1VVUPm
HmvU1H55Cl587RNiUi+PPDhZe+ETTCHDmAT023kEBiktaCSqPeEm73vNBZ7vYpId
PD92/UKjYbkKfwAbOHuUAMccYPrSvOZ8x4BYR2wQDiYrHMttVY9pZ2xAgSuqBEu6
XV860vmMx7n8qSO5NP0qwv1nqULvpaWngjRzRG2EdCwOCrcut4Xqjf/TRGTkTGsU
5da4noe1xjp8mDwShu9CKIKv12/vU12JkbmIFwCyitayLOSQiCU3ty55t10reS7a
g3GpfW7jvi3cB8ViaKKQfgg1WRHIiGHB4NI5C70ox2HD2FOEm45AkNF1gE9ETOUR
2S35D4SGLcOpQJGX67zPVAAQj77oXF6Hi2sFG40her3T89HLt/e3WHMQG0hIxuDa
Ly170yJbGR1wG/qozMrpLZ3MtMwKI9zn+OTtLHieAPAi9dNNKPk333SqEvax6xOM
2a1xMuD6fGVjYMAB9hgiDKmJ76fd78m6yGa/Cqt2gebeF/4rJZ1Mk+4q+Mh0p2lr
jreHOaOdVMy3OLBbAiajKnJ6qIPmZhRCOt28FjTHmr79DGwWNo6V7MTaKIG2HAXq
Oe9JUceim6rbLQucPWB3HPwMao9GYY0hg0luVIUFYGMXBY5y8mQMxSDTXqrMrJf0
N/W5XWXu+2bHxQr2I8VDFGw04eEWWjMye7/e/d9+Vrp9OOnSxMIQoxYOzrpnJXkS
/MvQWqzGz3QoCSaxLYl9fgYYi5oVfQADk8N1ggi3Tt+Qc87rqOCgKxgimjIixPab
Od1nWLrz9Zrr944vQZkzT+CgKccGyuy1pKA7DvyeUlDorcHKm4JnlOARAVPTIYSn
ko3s8nw8vduKtBmknOsjeuVXRLRDAdWsyidSEnW/1f6dTbHt7HgGMF6dPBCM3PFf
MSDOim8/VIu4WLH+UXwGSfKtzvMfhQUYkoL0cIG6n086mSZQfludMfoKDy6esFiS
U6yMTRU49vj1/y9sGe+9z8j69e2HpN/tx7lOQvUZxkanf131m8ry19/kcWipyHHL
sq/5n9WEV+Kago/fK9xkhLfxtqok9qGuIVbNJNHFeq/B5OZhf/DGavf3716q9X5F
VStOVHFlV8Ft3vpip6QfWqPNgpyoHHOxgxc5kUVk3c+AqtSBJIR/CIupxjpTQ/g1
m0w4iWt5tiiBEwo1oSfOTE9rY6YfCiEv9yLfU3iGeLQNsQwgHp3N3NAV/bIcgwAM
j+qHus9KAKn+r8uZSIP+frVstMuCeQhTPCt6sbn8cd6oYxwtQb9OFxS66/6AQSka
6hiSsaP1jSFnZ/t5KkgDPClfvZtDh/WC/Hk71mm+Y9MWOW6fRHCKFSeMK2ANvRXN
HYSowjO4AIEU/caXRtaTHRemyK3w7gnabaX6sDqc0NV7s49cLltPb0323gcvoriZ
AziMunKEqLVjAyQiYNN0lr8Bug9BwIpPH3b3RH71vIjOP/Ygm9qEoKYO9MpqAh16
11wL9mf3v8XVGJ9ntxk+J/rW1YU0QVdf129S28ENa0BavyrHQd9vovFMx3XRqN/q
TQuUobRayrijvcX2r3ilsvf/QFN5ymbK0OHhRh8WPySFYlTGaRPGPf3G0bjCT/Qm
aB2U594eJnXbsLSyFwVYXucUlaYl1BylbzLQwo4m6RDXtIsozaPk3Lf+hRmubDYu
R+pZbgc0kBVzGBnKQWE+n6NBH3ZIMdEPYHhutZj0FZEY80sM0z/jOwAE5CIU6RNs
vabor/rpae3TuIxXMZ1+jwPR6NsYZrCHCw/6fR4ayIwtnZ8pk5KL1Gz4h2uDtRCA
/JOtYHNT2bTEjmvJn3M7+/8t9zOwZARxlZrma2colvTHxns2igervlg1mnTlTd5+
pS1Z1zSh6bpn3GqfA34AAC6dG9QkejxG1GLF+CkeJ1/LCg8krvkTb+6qHcdsVh2R
50uX0gIRUqefMkF/HgYMkuDVN62E4KxFJaBGOhAycAzCh6e3zs3iG8KyrGOnDT5O
RDpsR8LITbh6UeRHBTl01MXFwGq27uFv2+C22jB+zkbzMlM2OvRvG8pVDcQBLwpj
XNRxik+q5z7lel+LIzsmEwIkZZbqRSAkCxYLMgF8lmx5HcaRzNQdEoc4LmiGc5Dx
FAKrz3nx7IUAGIaiiOUTLEQ3frFJlJq9k6LIooZ+adgq7gsDex3k+j2jOUooHx19
36J0p3k7OReWNZq8l0COU5sgeqAQ1MCf5Iue77cHwALy2CG1BcSN5KMr7Y9anwSJ
jVQXy3obAyJS7yCcigvyZLU9r4Puw+E6afFAyL96u98LgtI/kjyJiVuIFJc9GlYp
T8hcMGQ3cphcNaxm94urqJGuFfNTkQjaEI3qNU95v9E69esNOIltM2AGhUZSnYTq
ZHLnG0O68TcRjBOR9bdqz0FrSY+KFFgnHzl2bUxkP2JUJBcwcDhlQj+5SRWmQzOs
lwD8GUqJz8+oOrFxcpisY9YUk6cHQ6YgjBhQha2fL6cVVPQzi7RmceBeKb1l+Xte
XZ3kA+HYr8t39nype1RS6h9Ln4v1HuqWs7TQP05l20Rdgjvx9/LcLxCtT9PeWqqY
G5SDmjkOI3w3Vn5Yl7KypKY4yvlPfTs2RerruGwPVWYI5HyUYf/bIRxIoabyWEAb
NPjjHtzT9dMP+Q6i3qrhuVD32w5BPdOjxtFHKu0iVC8JoU0Z4FwpWlhyVaf70dX7
2d79YJBwRbbYJj/QuNz868FblN4gaitvIv8m2bT5jQ5TGbfvVckr2QjTgZhLY3kW
tcaKhiReuuaRobeIKvdKcViQ7eqgSeAgv8rObMzq6a4WuDLWlbgZCFyTwbPH14KC
0K3xYuvt30prrg6RdVbK4NKVc0c7s/epRoo06+dyniBtUendyJ+7oanirrJtFg2D
s2HfLIbv1sD+3u+TasCjb0bI6pnCF3HSo74yM7TVuGt5xN9dgtSTx/xDGYvxr21w
uNafcTM8CR8vZLmRjnr/cbzg8Asafz2eZmIdP0IgkW9OKpbKubAvd1IkO8zhWb+4
3oREEhEksyOmAfzmyk6MjYayj9LTRANzDSiOI7se/JW/t/zynKjtQ9bQMYYBy4ym
O059mlek5TS8S8fmxfydj6F81O22uyeWWBLNFBFstOOvx3kTROwSjfd+9+o7Z8ug
rxZrKEq9bSxOR73pRlLhIZgWlyWs9iAEPJkTOObdMRgZcZqTU/aL/7hUIMI2IOI9
z2vL3FUlR9w7UdkU2rYAZm9N/9F+9m3EyK+lZQm1GFm8XOJGGgsSg3VydJd3X4dL
Wmjf0vqVQpBMZgSiiy2jWpC98sbPXpPgkAfgLpGFpZdvpWcL+IgG7VVczfTa22Wy
+6J+F7w5XSHUiAHtP8MUfOaA0R+UWAEz+KQ79LJZFlkiQbgejAL8eSnbSjbhICgs
1TUOQ1Smpooqjn+Z1YJlC7BC7LsbUykWLPXLzmYtNSA3jDqwzG1yJI1Z+KACkmkN
3QKdqOlzreUQB8XT/9/LiMNT9jx7lK8sCya0NmsLR2lfTJnUf2a5bC7EQktDCpsE
8+XC1iPFMyUYeJ+iPJ5Ft91V1nxMjMIixZiQQuml5+yNRuRv9pi7tq1tz4tOBv63
ZaHPUF9jhaZrl/ZLzAvgcxb0p2Q/YJxD7K3OXrumg02YUuQrKeqjF7Z89RZo4uzS
xihU7C0KPdSz5YU5t+mgtnE1QmFvedEHwR4fevSJJZsNiilwqAGQOPeB9W5PM9cX
P8EH73b4lpOAgQFFDvdRfvtRI0PvFSrj5JrekfoIRdWH60cYEAQCQQbFeBN1+M55
A9MO2bgRmYuDio/igmv3i1SPTFdcHR0iP7pTNK/bSt/t7iZLsIWef+9BolaOjzZC
k3MEpgrFU8mTR/ymMXMzVoUlqNrZv/fTTzo+BFmvoL61WX/AUX5/2+t82PwBYuLZ
5YcW++9XZ9AcHU9kf9/5Xsnrd8jbiR3ovKckc+sEbiZwU1Cu4BXEgKpEPLQ0vZr2
AURYmtLp4Ot48hEOG8SIBD/O7Vy16yUl2xaANIvGRpQS6fTVvPMbGoaWtEGdYD09
UG9NaNn0oLz7em5uCYDSjUCMpTBJBJnZ2No9yfFRjCVH63eXGXh9o7ZWL4IU7V+w
nXAVo2Ok7/qyeYiyZ08/Wvzv65jd+8rj5pB6syVwipGMZu3buX1R4nHTk8c9YEvD
g6pihG3WLxX7jfdj4KYv2wk65Iclu1Kcj1BvY4Y+AwtUAbvbNdm9J7PIs04aHNMP
Cv3P+OqJT8G5c6apUUlfYOZhfpRAfr7Q2zejOjKFM1vtFJAitk5wvPER3fHHdHZZ
Hu7nDlBP8qf7owbW3mXmU+pFf1c4PafwbpHI8yWf7PcNEbXbuVTxfu0Pt6Deh67C
y0CfDpdZ4xnjnJzqyUw399TOaQipNvcxezBlyE6J3mtrLUCSxyk7m2WeeXf3Snw0
yybV4+PTsfpc26bFAdqqGws62L3SHC1KUxN8y2E8oow9c22Yw4hTc9BnREa1kOxk
4VO/FOijoL6N5SzLH5qcNkuPCnWgTbmHkgdja09G7s1uX2IIDqsqda/Z4UQeOVwQ
v/CMraOF+YxQ6ffo7N88GnCXjVt5gqTkfA2SvkLDHy8UXGkfKS1G3viKw/Qr2EEi
QB+M8ohRle14U/lzTjDz5BzLl0aqrkAK1NVrSrzdFWd3e+gHJIxCOL2BH9YRf3VJ
f8sU+pTAzasYTU2DDajeaPnEtfs6M0T3m3JU1m6K35auaj+XI75cCDcaYFFW/zrG
VwcB12ya27zTJ8I+KZTdm2uIjv8TUrfiTUyBIk48SJKUrhhzxzgkZVw8oyqQ3IAy
OFS3Q5UvJQBGebgu32hhHelnUqAKrgF4T8KkI9oib1cEaoP2Lel1m2gH4H3GhHlD
zY6ZHvgJ5uOibBshRVV3JngCF1McogZPy8IGta9ioCX/MV1k+fN/sQce6PiegTKm
UuiCtd1RDSjx7Jdq/jXmvqh0Zyhcq/PFcwzzmnBf9WT7qPaqAqLa/ayIYaolkSaG
XjlPh5wxRuIAOnCm3pwsX5QZwPdsY3UwZft8mE7ZlPXaiF0vkw5yNMSOBxvQDVAI
Q6HB+VmiYUrFp4PCM/vfBZjGyWHo1Zu9GJ9ZCClJAQvQibByrou/m5wiWC7uixiT
cfk+dV6a5mAWKScsdLcDBwrKjPI9dFLGVZ2GRyGZcEDzMNb8g9cs3JRufznZngMl
kWBQNY5FzbU2v6bfN34i2WT0cQE6gX5Lv5zIRSVHUPkvr9lCMQKE/WlvTuYYc56u
C9TAyvbwRM46KjmdCoqMEsWMCT1S8/tlK1XG4gZJvJiKPjNv9Wpff0lSCQYaZBg1
jlMrnpKgLFrG+DRTJFYXLDAAJYAHkjJvmkY/D8xi+wy3VwtKeXfmgNAuCT9KNa3/
vbIJzQA2OYULK9LcFLUg3csOO5ermBAMI3MlCtZmAC8xbXO3U/0KeT3B17qGNSiM
0KRgSkKeH7KtoL6Kf7gzcwkqKAQ30eSpie7EH+torZ7DZ7/9qAS4DNcFfmYVpbZk
jOdZTmUHuNRyjCPB9/5EDjcmb0EfwirtoyDIGwt1854ejn+sDRL+sr27hgNsnsLr
ZOtEvJLJz0JGBwROlqEL1SnMRnU4ELC3jbtUtJJgGyYSXwvVtZC6yev8QQT4zmnf
940rsaKOTX/oOuFZSqdN4MUAM201WKYM+eD5sOo5YSDLToBBylyW9PQkKyhdL3Oa
JWg6kkpJN1bE0n9XXh//6Rnre9rAXQ1E6LYe3UVeOt+Jwvw3Q7VSl2Q0Yzj3vYzX
woQWhV04TUnIASRWEA7qPYIcV9BlWj8N4Cold5yn20cp/bF2MPeJansLAnLWQ29E
1ehI++I5h8/ojZQ64316p13qsQnIceq8DPP6MG7TLrqxMc/81Ijo+x6K5mr1yKoV
qIveRQ2YSHMfYyGc3cjqbvQHtss/zNaTO28McC/9GgaGxo24ZISUTUxzocFDbohu
EMHFOXf1jnBn08K6HFnSI76nbTDm1CD+rU9fGzI0sOmEjaaMqyrL9m/0Y7hAZc+w
E34dYBeoWjihoFnnV7Zbu3/b7+wVVmxVokRYP4UxpedFeASsRfdPTUKXKOa5+Ftd
jSZALhPhHWgphk48gd4PYnNtm9TeXwFObpT3EGg7lBFlWYrRgFX4/0ujwT71i0cy
ZJTBRY6Yd7c93M9qX7G46tZcvIaQD+c5vRymwUAqH6L90tawmHrYH4OViLTkn2Vs
StjcFlIaN+CZugSk5YbAr5tbyvt1SbstvOpExMYPUMEdNS9Beh7fHkLb0onGaUpJ
BNv9jRWUr7haGVBnDXKbbncyjF2W8m35WNZPXkXh1C7hQCOF9VA5zeGG9ztaI0wY
tMudMGG1/oUKf1XSEmMdKzA8yacrIrLxZnQKhz4+nqLuQPJ+6Gwx9vE+SeJoe5Rg
UVOp7AXfMfTLXEsr9iU08U7s8QmYiF8sA+kGVc4PsWq70Fxdg30NDTxlYrLa9HPV
DErxWAok7B/p2vM6o7khyvr/ihFOggihouW7mVn6Die2qnXHOSv0q39V8UhvqXql
irRqhyEZstIj6FEJN/8dDgriPkcYWI8OKKv5MI3JMTiyq0bXX5SFDQCPQZRVHCKh
2xQSySLsYKtinJwa/3ZIT1JKkAN41N/5ulJpMVi+iPFdzAOq7jkqPhyWUMg90FGX
ba3p+qUNQ5IbO4fWl/oHF/rgBqG+PSAmZ5EBuyt+aiDnbdFKtxqm7no0AK7taRgx
CA0zEwOiGNnJU9BVvsveKcYs9ZQtqinEhPhHz6uFexX9QBDfQ254Ed7mk982GEXj
42BqqkKXT9hQNxNYxKd+Uk2faHghg8e0kwUYo+WYDnXxDNjVag82BoMijwFzh7VS
xOQi1VUx+0Nxgy4UoZ2Do3ouFyRDQTpsmDxm0q6mxRCkYiJzqOMdBKYFGDxTLGNG
dC6Es1TP/K85qxCVlvkhI/zHagy7JIgVu2R0qCJWa7XwPDu+D9pEH+1/DoIRCMAw
pAnSqlBITqmg91W27JX7QgE/Q9ojiOad0IFbrTBYBsZfcT814PhwHdUYH/kSWY8M
3OWC615cYygUrGtzKfCbwJU4ueBzhObES1cV4T+0dQIVR3VGRV4iM164UcWmaHTa
jkoRJOPB3H9PD88KFBS0TWqUyqxZT50ijp7RJt4dnxKwj96g3PLmNwMEvSyl63lC
+LpOr7Vs+a55mkKR4Nk4AD5aWaWI4vjvWfVpmsOWNMcDRtO4eK8tqGB/PXr6wHGL
KLTSEUh30IpESDufZx0yMXdR+Mu3sU7TTkE9p/W0lFV5fQ41D9kfkvZE7je6hrSl
1vfJ20wpgofditQ/cW5I97DtkibX+FwR4oSuAoPSK2P6vB0AUAIYIn2DANbAzy6u
7X1lPZ/5YTgEPtFENMH/2F55q1JKYvkRQeZTnCysMTgQeoaY7xZ+/fkxMxJeDjK5
85kFtax01LvDG03ZhjHPYHqA0/2yIq/2EWAucGbguLQWxNlVWO3FwItnqlmk7he5
6ZVWdsyLi71fEsnNNLhxywKHlMGYLhOrr0zs+ohXxOJoVCn3dju/HFUCmPCfrs57
kIrob/jsujfHRDkRfKrF7w0K2kfgnRHVkK133Izfr6gu6E2tJ7zsguMmvbsw2AZ+
qV6ND7Xo8SW3QzDEtqHiFSWZqzIxaPUVVufY2nMAGUyKTA/KS9xu2pBw1a+LYg3K
UsYNtJvwwi7/Asw04t1AzAe6jD0uoi+6NNPxpq6w3J+7f/cx1af4l6G0/qCtEISN
I8Rapy+28Drn2TXgGvVqJ1cJ8OhOK1mihFi6FC6QM5i8ut5e5olavG2loOPCcuwE
Z6yKFwcz8pNgUXldg1WUmMFXTGfohQlhlwCHtmn+Zy5LW/xUViLzgSq9bPbUbF6k
XHw88wICr/UYcZLeNk5MpoNF1FpOoSrrYm9/yfdOtVv/tbzjCnNJhx2GbT433B07
MqyzNzYMUu/JBC4np6i/9wrQBL+gjScriq/uVuTA5o0C9EMeuh7UIpsEADXc20fr
0rpWyRv2Du93qldbGn+nPp33vIwqWvG9AnJz55mpJQmUKtm75ZBMsJJQlhKNqUqy
KDYGXnhHzdTe0/LHVXnrvVGX4l137zHk1bkzwAJYh4B34Iru+H43ljIq/g7VT6U7
N9t9ipXssw7gwytSnETp6hTkFYXKBi0KrmMM9b7J8N7nU7h6buuKe1600RZ/0qRi
2EZJ2J0BpDNFOs877nidmI55htvA/ZQhc+YHgmlYbRTdiPoimDnBeBlyDNyiNwIv
G694nzGSoglvcba3v1zVdALtZKK1URd+W2tsk9XDODWw9vNkGi9vU8pKMSSO7XrZ
5t8IifsvhYToe5buIwjgSEvd4YLbVzoLvKPdpadYVAixMFlR/mJjh/f3Hz8vwMvz
Fsr+KqAkI2iOurOP0qgp+NgcjnBWG7zVXjdpICIvggquU6w0DbDO8W1k1f8ZbE+U
PY8gdtovA1jYqqcR/oWoVAtKe5bDZHXykY2hqNqOLVzw1yyFOqv8SBwvNVfNe0fx
9qYJ1Vzl+L6PH0pYUTs1kdhaZNUnEniFNfkSZj89Y7jHSN0B9gy1alP/nL17YdNK
E+/+sdBCRdH7Eda5aF181j1lbor0MXWUJKa7OfT0PFh/iDKIvtuLztW1dkwwGU6Y
t4VgO5YIz+KG8CRvkHurBu7zXGvhF9cagqkHTdT21/0v2q8XSq74iXCJzO68Tpin
WrgPBBmOR3E0rFwvo/FBgSMEYyAP38ZUJ3s+fD/05wSBqg0aVSckzF5etlCWNHut
NVi3FgEF1tTqsi9fRm+CmBDozXsa1bLWicX8l0DU9tA8GtngMTTtKGk9ben7LYTm
90b/hyce8TIpWarAv8js1tuREINo2V3DdhmXOl32KNhtMm7/l4L/WTUd3C7UkOKa
Frvte4W1DMomnBt0byYmFexF8xz8yETwEDbuYHJ0u54Zxx5FCdGYY8VUzPOkcihN
CoAvRYH3hqwYEvTfHfse7k+hXb/6Gw19dlbZXiacKuBZWU3VxFGhLAXJw1YDBTyR
SDE0lq1uN/8Xs43zDMRcLILoOxHQFk0dSn88Oe/zWStCQasuU8uZyMLOcoknJnAh
9nJkhdTwKDRFuPw+tBr/LFnW6ANfgTR5gvPpU9+to/4TM5Si+Z3qlX6vzt55YXIj
aLNl83EPt/7hWB2fBiL0nKIkmzgmSf7KV+cgHUhv3OWkzv0rYO2bk3tOOzLoSFyz
8w/NHpfC9MKMzTJUY0F/ktEpXiZVBHzVjw11R/DvZ22JVwT26T4MiLhaIPrePRuN
cZvjgiDL3F94b7PQOUH4r+JfczX8R3q3NfGGZCmv4mY8806kgO1I4MaJdjLCiQ5n
202kIKXoI8jNqenzWphMAsaO28mtLOgmKJ3OI9Pzm3fxF4QorTdfdXndyJLq9R3v
U3ophH8qWSBzFHvUnut1eAHjW5Z9+8Wh0MZy54vMrHHjGq99ZM2jBx24UI10EYJY
8xgUapVaXMPSFGC71q5z+By2RR1nhv9lqRKxCszYIw/fyLnIVpd88WtgUrNghge0
mSF+gz0oTc1fN3YiNLzJsCUeWlTOM+yUIV9GB+vHolGBR2JQ0bDb+JkGBIwmaIWH
3UZNlnDw6ZlQlqRJklun+pl3V6a6ZJkdiPB01yDnlpj6mj26dPuKEp/k8kNh3oq6
IZ4/Zz9H3ssRcfXw7++98ED8r/r85QuKbGzvirREiiiztuhmnURGfHFSciFQw5zV
t43iEAePmYPHY1SCSCOEIFku4NV2UnF12vTroOQuaze4UMRbbkW4gNl2P6tUpjW6
3TAdWiYMBmDQr86v2AP1j9J0/UrITDMWwvdZYChvxxiDEPYJ6d3zDC8C1IdjEkws
ISE+S9VpHzVmsf0OBYk+55wKqVdqQvpx+iQOzAcQJUHoG+WU5+m/gn39Lsrf6Db/
UaKYWS+f6UB3Z8M5cHKyGHp1RA5T0flEdD/C+xbsu9ympy1S9Gsa0AdMaUVoql+l
NgSmRRWGgxGPISjUjpop8Oibpx4u2l+pkqSDcXVomhchYrCtUsvJ0Ew/CBbJTcds
sWcUU/qhiZ0/9KEmQxrxJGCvReDa+eePWyzcjFqIepCG1hsoZEgOAdNTlegBrwy8
OvZjJ4Uuu8/E2DM9/BLcRodzTdvYNyDOErHPxtsJiSXHPYPjbgwvF+aJfjm4EIW+
a0qcao4BcW2GQX5n76/FFRPgBGHHWg9lIutMX7IlWJLwL+s8OY7AMbIPQyED1otW
dLTZ3SQDRzuTF39OakZBJyydcv5HbhfQPJevPev8anfdoeEwyZupTuqP8TxVSkEr
B3HDPkZddDL2+RWuc3Iy0fwv9bxBwgNqvJdxNpvnmo9SM5Gjld6P1+EDnbq+njbL
IlRGGHJOWREYvV3ji6J68lS1ELJ9eM1tCv3YdXiHFggWtoDH1+OdX4mBB9ue5xR+
/6KjXEoJ0p8iNvBlWJJ/7b3nfEw1jSUlDiCn7ODee9VG5qbM95H+jOkDECmbI3t0
L8ERbQyJ6g9tNfao0FwTq3ToqntOjywx0HgvbQVMeHWwmXKfqfoHQRxLDr0WCJoS
+78mPkP0K9vuhAZ9mKe9oCLJfxlpv6kMSJCbc95dYRLPL2X2hqoA6xUMSMVJwfRc
ixpwlvQq0lIHxxhBXsk618BnynMVsRLzXWEyQchVJ+Thof4nCZKjm1ztev/NeZRE
BORYg1IEfXC/Tww51R1uW/x5I93JWOgPDZS5gR2CyU2gecu8mRNuwf6lIkhXb8in
aHaRE1YI7SXPnW+1aXASfsaV34xm2NQzrJi5aF8rMEhrPKCvlz1W2K2ZiDE85tCA
X9hg1ZbQfpVZ4rcqbyljlO9XaRsGo65+N108yNyrEyKw9u4uWRNaY30aYSUxBWKO
WnaJiNVcIPO4iZdeRLb9zc6K28j7ZHRAo9RhpLp/ge0HEPTRPV5UOoh8IGsX015H
qpdnKI1kPH2gM7bHtfRa9M62Xc0Wc0Zt9mDxaDBlVCv0fwQkj+vOSNOlDvMtPq56
42T+Xp/L0LaPSSrgQ8n6Cr9ReTiTsUcZnVu4ax5AZNiUxH0U9rUIUWJ1AqJzg+Ph
uxpAZcJoDF4oRDRKQ4FymJfUYE12c5b2Lk03w0C0ehrvDMUZC+J2avmFezcKTCWD
n678Y8T3c/SVF+tNVAWRecsLHPawjJerudPjqhjs7evruEjH15u0i2jI9mqtanA/
qcFghp3sjka9w+AGpgJONG/8MoDvbuXed9Hw2Iuv4ooIZJiPpuuTA8v7yczJ1vnF
Z8FPwl1FStTukHlD3vp1FW+siuNTlHwSS9LjN9uHDDHRbwBaP6FVmnMAcnEqnqIO
ux1EtAs2aR6EwOY1HtY8bM0WZSonJ1XMrQ8QZrVTudVF4yiz0UKQjYQwz9UeBkYW
Mqj+rWKjzrbIkbBsAvOtZSbxmiiuqMlASsJeGiTmI+9w3jD0dsw4z4jbRNCd084Z
KXThdnOOEpDPLBz2FtPR8KG+C9Eh+IFv7s1VWw4z1SF43ln4qPNjZ0GBRgbSAfIA
NrviuC+JkZ67JSExRbdlCbIIst3aWrwnLTef3UWFCH6ICgpGppPb0/bCxp3/puPr
RgM5ooujCkL2OwBIsQQdoUlznUrSG1AFpfJQO7FdHuPAajwjz9EvdzUyID1jIuTE
NXoLZdbAKHhlL16aZARTLdu9sg8lLBPxPDMvurIBjmIkVjrJpK5HXHyE4v1hWh+1
Gt0mNIn2xewq2+KKnRq53jE68YxdZUbExXRr2m7GU+AwMteSjaA263ccw6+y/R5E
NI+dc2r4SR5sqogallRcVtTQusgyBkJC4o+MM90dXB0kMUE7zKa4U/h1loE/yUT4
sKyQA4NVfdcAuNVGJBO6r82HicgAxHMMpUvPL7C9boflZm2t36Gu/9sb+BHDDwFQ
QZ3ztrIzn5zyicZemLV1mcgPJV4GMoxgQk5aGVZzQxkf/u9aRmV8rlOaj3J7XLo7
GtRACfT7daL46/UgQKykoQxQUNBDE/hbm7TDJz3NBbUCiVqtoUdxPnwQN25wqemQ
J0U3TIoQPQRpKFLs6+/vx+tJwqTTDQRdvtKKz9kLfhekjn7MVbUUclPDVbE1uPL6
c2f59sSurAoia8ImERY9yNkxJ1maqFZLOf41crUXG8GuzWWJhmYtLp8GyJRnMywO
ylECKpMKe53fEESBDPK3mTiXuCMKhg3DkqzFtU8casEnNyKu4pnzs1SDQ4sLR6q/
5/LY8KOsGxpTUhQ0p/zre+rfxX50/4QQ7EXgNBX2AFgXfNqayf3hX58I2v5+uFQk
yvw5GclnKo2HnOcPZyDr63cI2nAKzyffsZtogkIl8zdUUFhEfld85h5fCxPdK4D+
9JmGCumx8a/8y6rXsrLNYjY/Ck85SQei5TsVcu6d1yjlAxs4Y7hF9ru9ZCBGy7GF
tZq9y8DK9C8fHXwwLZQUm+4DvR/cgbOr1AUAw40B4QxCdSO1Sbq+kBjYi33sNUEQ
CH64Pa+LV0oYiTH2CE+2vcFRz9uNBVlRN1DsLsgGCfxIo6/y4KI0HBy2DDPgFg6w
+3e0Yq62cI/tZdOWUR/+ogfYdC1NqRwm2SsqfMtWLdX0ivR0Y6zzbg8qYtBTQuTe
YB3Vkf7kXwTpYaarSjM5u1C6g6WhiMSOd+yeIQqy4Yylu1/b9rfVaOlMqtsvZqNW
jRvu33C+eYuB3XAOyQ+e0q+3YpNOhMDtEZJRjSjCPwAPVm515g7MxWvYYy+vq21K
lYAQi2M8jlYz6sMcllCTFkeNc8e5v85XW/OXrNNJDAZsz1qwxXhqtXVp/Esf/moZ
Vkev7UNQLJSz5h2TEZEWDdggF09G8hXbZz0BIB98JYjrsgnrrghaR5OVBTcYQPuV
QxGSFbhFwLYReQTOFn5n1kTgn315K+Bi8clEpwMdReKolySJPoYecJU7aYz/8Ig1
JGcUFUltpTT2UKp3DKDDpiaHAe0xxZ1jCaGEgtLFm86EppIFHwcrx9rsGmEpZcY4
eL5TtrpTIFy+uKW7oDsJE+BPKFfA7TSkPsm6FJmUcYvwpYFb4/UDZ7RjlCFTOtuS
NEpMEbX96aHAj9X2/tlMiEkBJjnneRlKPHbSDVhgjaABPi6i2AOm4uXyCJsCo4Rz
7fn0OUfspXAnSkfavsZrooIWGYdV40Yz6NoitHifjaVN1SxGldbUtQtzrBIjsa1H
prM4wma4ocPl97a4A6XUSJJrcysls5FPS1Pr+58MpZAJ+P7vdMKDaUTmsN6tVAJw
ygKEEgFuhhddZAa5j8NGfcEh1Xg5RmQpa0kFNzBJPn33LkkOz9lxOSwQ38TqDU34
KyuiBV6UEX9oUBLJPG/bVxJAsfoEWFMeqdgAHBVgtIuQws/zGRkKQYx8rO34DPGq
4dA4sxX8tEhGX/eFKIxqFaDrI1HsXNHgZrBes4Wax8OXBgUkVzWTOjfY2uV6YxbI
4PB4mK03f1vgVg8ilQK7JD8ATW5ZL0D1Jy1WLp9MckLmw4MtCFUpmVdlwYR3n+Zr
Pv2+ucGkQVdDGGceKGmI7defnUAZgWuVCQk7AuE9RN+DSk05cV1GenS4efwIepxD
2P4L0KjZjc4GsmiJxbQJCKBu6q7W346fzH4jHoTCk7Cf9kxwY2onU/pSLptGfjoT
PBl9gzMZwf7oGD/wHIcFKAKQ3iAFKZeYoDlvxore1B2QlXK1e0/w3zPLw1PSQn5R
Sa0FsMUjEV3WHMudepPZ7kXp6V658DJYRtOzoWzE9XD5kZ9yLeDPuPawq+jk1tKB
Mtboe39wCLvSae9BCm9dDdXDtc+ddoQD8p4ysPibKi4HRQPZbCerzfsxIKcw7yNV
kvA2KMq1aEqrccXCl0bnvonEhEmB2dBgz8PVk+MtKWEqkh9ezz4QYuUJahjWguL4
lJZIvNBd8MeGyMjxm2Y6InVJMQPYprLhshZV46jsNraWMIhp6pAM+XTY/sAYGFAs
EowVgTVnvfhjjA2RK4ZIk527UzKayq+ZjWHc6jNEXLDhYWj0Kfdwpa9HIembQf1y
6/EhE6wZgZjJJm/yRV68phcLO4TLwZYVFxD+eZyW9mD2LyJmwqPlwnrYObKVMxWQ
TXBWcIWYszH4JtRmbY7RkYW0RzVKm2+xs282AcQkyHfOYACSFcVWORuELJIAAU+B
h2lJ9Qpn1gkZgAbtbISSwAp16HkTDbTUsLreJWptzBoeSOkyoLxPEyw0NSNhaQtO
7hXqoVqwm0fZaYajCn9TttFBkKogdYEbPsIZwZDfZUYmX6+snXUzkz6jNqeWUrG/
+DnOSXGKEU1GqgCo0gAo1eNqcYxeRHIETKMy5VBrr6LX9JjXJavcMH6OO6S4QJtg
o3a70/g50OKRSAD07H70DUDl1X5YrEvbM5hPgBTMuFMoi2OwxzP7Lbfjrr+CJRat
q1+oJXpTbGyH2xZYwgO/NJUiONpPih7Ehi5cxOfmY/3QiNahNY8+HbpNQssoshRa
ySLPZaJSASbWgTXPZL74nl8Zp8+3HvoD/2evN9DJzJ8wPrcS+aaz2Qf8VHIo34Y2
bmu6KdAMVGwyQPaYbBjGFAATiff9CJQboYvK85rh2dT+PA6mOVyZY2m3qB8JgDmU
9te4JkyOU+7lgVrf8bAwgh89Ky/4E1QpDkT0+di1cwkJes8d/Aug0aM3lO11JCyL
NUanBWhI9j1AwS2Dht75igDyxD9PdjzyjKVMKDNiUQM8QmFvdQZU7tJOC5iX3eKg
4IIOjGww4DvXtC6kjXRu24d5xv8rODsC8ImanhrhtLpq9+ohCDsNFKRi7eLhH6S/
81FCi0diC3QfRac3N7nxas2U1tSfvmmTUiy0UhPTWytGLml7l5j9K/w+YPYcVI3T
fZyODr7Fq6NLUdk1bOm6tMtwb330SjCZLQp9VsEgY3tBqYFOMveLDg/rXyxwtGZ2
2m1llUp/fGNVl8YRtBm9RlT4VM9kfxcmDhiMsTBZ1hrF5x3KWglyEWOdH8yEnxUp
wA1guGXcYU6+4aaz6gWmHfp360ZzvX5qZ80ElGIw8qpPpefCh5mjxQERvQezjSIC
z39TRsS+gLr7WuqiZKfogOMmSltOBMU97odpN9BC7vRzc2UKFlEmEbYuRmLzBCMs
fPMKt35Gf4VWenuAGeygjs4r3a9TiwrZ+tq69iD9pfjutXdInlh/25DtfSRlfOCo
2kC47RGkc5rJEk011+B5mz3BIKgxIMShnU7fN6AcX7qG8Yezp2zV4JSevY/p9wbV
jCfj84EEg8ab6Wwzhtkm6J0maeYk2XTv6j9rr9H5YK5kKOQNN+FZSbaYSxUdp/wU
DmDZP11QWQFZCD5Db3C8Epx8jQ9e9+bpD5eJmwdsPk/DYWqaFLRV8FZ2RPE2di9q
yQGR6LcZX1lsg0rwIv+cOK/I7C+HfABWcf0u+uSYd8dg7oyIHvZTrz2kALqn+2Hk
BtclNN16NnXUAZPJWd6AHfp6X0xOTTCsIz8LUhjgVi+5sRom9r45KvbVUscb0xoi
n6EQwy3uSaIi2fM/pEwYE7mp1fG8LL/N49sJhiunRTP4H460gMnpsbmr+EToIApQ
C74nbzKgvxqNPHdf0c8tGWjNK/I4he22mjr0zIQBPeyrGdILn7oehP01SnpmP0+2
e65/ZyChc/zu6dfE7u11yfR6gfK5yETSM4f8n0uPIAfGOE6Zj5rt2KkEjH1pRfwV
ytM6nFoM/epAz0FKMzieZFWlRFvs7Zwb7H6kY/Eud1FXg8bw25M8sLH0pbaKm8mx
GjxT+AUBzjIDwSXf5qL9LMwEhISqwJlIPTedHbwYVMyyiGlJ0nfZigReAwS/HNny
VE5VQ+vhWZwqsPrWaNW6mRo0GcLt8ZPzJdHtrLoJrgmcCIbwZn8nxHAKU1dR3xgX
A/dZcbdsp5BxMcp/7wYGbQ5oa78H9UNX+bRik9pY/wbkVLQfTOhC57ZvyL+UvAk6
F+zkzpLErVbllQd/jGZOSdIs4eoMITr+dBA7o5fYdi7NH1ozO1LbjRjB0AofWzPR
apLl1lpndmZY5qcob2+y74Hm7b1xFxHITBKrvFReJ5PYb6i4ijnPp1/ec7P9GjvV
H/Vc7W4tNQ1t4WCQemP0YYrYmOiiZXTuWc5WKCmixUJlKG3drUYeooJ2rRdatyE5
AhXZqkcYXKM0Z56Gr/2VPu4GhJJ+wiQaZBq48j9+IDcnBSYTqRKIVCuEFXrIa2FU
Se+99jEMD2JvzeXczMsmphyqHTKpiHpUtKAy7FsUg8+efGFXZU3k7xBWNrO25Dsl
PSYmE7r9R9E+rDRgpROod71ypE+bYRCtfc/VrZVN6sCM98B54FjS+HotnhkLkF/r
/R4QYGQuHlwt4OYvbky904R5syQcqeM250ifzU7s5qDHiurKpOiowMokFjzOmNsu
FnRvwkACyGf7Cdn6gZzN/ZeG/du1L2lcaj3fxZrDzQWH9rWGMQdetEUjEErMgclL
cROJzuwZ7sROtJLviUh7P5yYXf1rSVZPDoGl80JHoNN35SSzx0klSq5yYDj5qWxK
vQBDxzQJFSEjM41Znn8g+MYntJWZRPnnq8Kl/pm2fKaZ69BQDhLsSS/5Rm5Zc8tw
UPiOgiVkdPqoZA4q6ksM8TzqV/nBPjMsMuRof8y1hQ/Nu1n2X/3X2rDij6JeysOr
dXG9h9QK4g1tXGfJw1Ozksd7Tr0kjYNXI+mqs/8/QO2huX3EloGJHfqcDufCeRLw
EDKxMeCLgj5NNQBKPba7EUfNPW7+OA9uhdGx22OMDeT6a27zwps42AMVnxUI7ABc
RuNVHDz8A5jUTq3G6Wr3TwNpi025dzz67zG4Gpe9KnwkfVUTDhBLVG+ivZ9PuE69
rITpERpWmkwbsaYx5ZJH2jXLFy+Joyqe/P/sGdVV2XzZnBP+1V9B7YXlCBWOpwYk
klQG6IvtVFosd1secyRoTDHOB8jtco8BW/+yjKYM6z2FDMM+ci7El/Y1Go+Zvdw1
VBIit0+lCukGbP8pUl6AZJO03pWX7mV/cIPymCvJZskxXMPNsiiklTMiGs4bk0i2
DAgG9Er62jUTdq6JpPO1oTVLXlyeCne1wowB/m7o5w/Cr8rTQKrcOjDYxpDWdnZp
v2rv/uupaM5J+E0nBPQfIvA4BaYlRkGM5snP+U3fKrURXqQV2sIQUTMR+qZTvOmg
KushaDhdYgqXdmeeHdfhtTD2ZJR62RYG/VyWfjzkyX06Gx9tTsdPRaxH9tsIaeMK
TBClrU13QRykzI+QtFd+UQabpmvh8H+0X13/kN/zTjTEHnbLuGfgKpN+VWDQ4XMm
qp5//uWzMbl5PyqZfKh4bmBbkVzF+zvCaji0TbtZ9EPD+REvMwARmB/k/ccln3rj
Mz9weez0zmdxXE8Lu/sCJ7rmHAchJQYiFLQIFQCqkUvuxiJgKkMODg8XObbm7/Y8
q8OS+Sh+eatbPxrlo3hqJSIqEp4SD7kpS9qdDsY3eHyUACqTV3i0ziAF5s9XCKM7
T0UV+NtEqweWxokmNoVU1W0uPrZNNOpubiqltf8A2rwzaKYwK5qhbS073Ecwz265
vyJh8BavApeF5Nx8G0SJpgt8auUAfPbFDE3HRhEnrEUSMDHz36gdhn/uToYgX7Ut
fYlRdOE8as2xWLvUHv2CYTlPJlxaDD74ya3Ebe496SDXvjpXJR5rX2fGPCuQSpP2
FtZAuofiCA3qSzeoXAmHGP8Yha4Gq++j4d0Tf7vVwmLIG8fl50vaTwHD2rdQfwvf
2QQ30iGYV5aWYUH2GuBt1N8d5KH3Oczm6l2qLRL0PLXDrraJ40686656CQP8sS6b
p7BXHfLjyegoF3suCUZ+SdTdPkEFAmTbAe+Us0OrGHGj0cvYti+OfjRoWZLF1G76
8CK6Y7aMiMhGPqMEoduhvBFxBf+/TKPQzft72Je0T9wVr5OQlqIwDe2CmHiJn3kt
kG5zoEEq9EZXTWLd4/b0NCECLn9XkpyTUhw/VdNUk39Aun1KXTuQikF5akDPS6P+
ao6H0L4PT0ZSzgNpJ6Cy/+JmZMGgRGU9bXAgw1jiHtcZaV1jU3cKHxavJvDR2Bbq
NH2hscdIEsHTJD5V37a9XUeoIoo5a/XPIdJ4BPxk92/iPihG45w+c9fwwCaoz2dt
XPCfZaePy9BHb6DsMyfBkxVasVvZ0IwcmwEKF/HbN21lQVKPxSt7w6VWJ2nnWU01
/bMOV6+cA/7sBPfDCO5cZJogFk7CMxu5Zm9/OmXwfhDeO4bwwmchQUd0extyNsjJ
zp/krVBtZQl8fs9r8ZQZMeA5YbZuZlw/XkZH9YF4N+uaTFa7z+VkefHlCbPG5rf6
Fs+V7k6BBopkaLAbaWuPx19rotyHisJDYdUmnEmilwUhJ3CICiXuwASrpNF6gcGl
AmB59W3N3RxHyOc7Wl9B/lQYiIgePWblv8P8XNpyASpNSZq1qxRu6t3DB2LuDEEq
ZOM0rrOZpq4C4Sh4v8kqSybuZHmpNOHvfCrW7VYlNQyrFWtNPxthcOVukAShcOlW
RSaJ4HloyvnGjJ34oJhTOB0mfyOVG7ERJb1U6mGUCKmAnBV1Q83Ydg+8hQMhC/gE
SP2HNbU8QbNysHIoll1Gt6GFbU6d7CmDRjTjfL0oi9J9GE5R5ZsrH3AE2nJqGI1f
srUvlxyFcMza1MK4zpaBRVA8H6/fj0lKTSo94QwxZrJ6miz2c+FTdNmcVxk1mAxE
FTb/UFj+JnP99wT8d9JVQg0DKN2EpNjkUDT8H0KnShwcz261meFqve3naqXD4o9I
QbxNfsnLcg1RlH4mswkxADULfW5ql41UHi1FGar0t0uCSVKAChNKFSN546S97Pc3
rPwGLTAn31EXbhNdt89lmwKN0mAihNZIEtZc2yVrRIwfUkeirqliqY3fQZ46/g4c
Uop4FlYd86IHetUYXpfNgD5zSExZLXjQCBSLVJvBRf9KRSSzICBqAowsElWQAMjf
puzGpbIE8f1TlXZyhST/hvUhm/dw+KWSRElSIe60vWVisEjwLDtukt2Zwm8Js8Ex
nmrDPOTcyz7svqj/BfoJ1IUXukfySJP5/dm0F/elq8KtdM3mge6uf1vK8QRg/0Wo
Ab/xNRCOwt4RRIFaNkGswai8a4Befhz1POvUmHFohJczxbnUtC9S2nmIXsTTMfeu
NHH776YIz0RfwdeS6LRPmwE9BHhQLHpKXIsKcoJMPL/re5hBM8qDTuxZ0cI6UB9w
ub6xAJmbgbDHNM1g9HvsZ9uwfaUlpgTLNZektLVjTO9S1ygD9D1B4SfGePRVX7ob
aLnDt1VgQLvjy7KCkJsu213os8OYqv/L0MnfjYyV3JXu7pwD24aOiun/lenzvPYf
fhwQ0UtStKf9cPtEJ5OowPmZEkfnbneWO+gBSRivy54rkszTtAWPWritVl13AVd4
a0NrToLpXaqkF9CuxFDQRU29kjObn7agYoCQNhKacLGNRG6kKSvyJGb3oD+4o6gA
WY+V1vTLCpsx5KqnkoTRRLZSpOSpc3gougJ665elBKelOlRvDOvYiE6fAUBoFpuo
KaN6/JkQfxHt+kT+xHtSj8FslaXXjfK76ykzD5RpE18gDkgVVbCrHuHLneRsC4v2
FDcO7Bncsmtda8Ashj6pJiCaOee9CDDLWUHBhT8jJ4IajSW/bbGwj9lq1GH0aPK9
338BWevzIi22LbWjEZDwq7d1/0zoY0fjE/CNRxlYOIrT7ZlVa2jTeppJaIVk3Jw2
4ZWkBksDazyOvhHr1Qbab0D/U6D7Q0CTVhvOgmJ+0rVIsf1VCZ/EMJ9s8Mnya0vL
NoR4IUtEkCU+U0JV9DOEGbrV8rqWCX8bQ7d2A4YagEvSbcpRQlRPEUABprnfX9Qk
ElgMUmgsAH3oERI5N8bfxuPElhsRQBBBcd+ZOIzL6Ug95SfG9tgivh1LAMDRP740
EGXcudPup5yKC02tNmz3hhQ8Z1pgfcUfWFbEUG6pQCVKzxP+o61YivJ806/fL7ce
QXlGxZUSX5v8j0Y1qi6NKAJDIF967VoapfLlDv4zXTI8iD4sRlU+/GvCUBQ7DfNS
HTZuheaLC/EtuJljeCalZCaqfbZYb3JxNH2ASbiC0z1DHy082otCUwvwjdeiunBN
c3hzRu+NLc+QfirhxJJeaI8n6vNwT5b99NkLMMurW1PLtYVYk7MceLNFBay/8cja
2mbgaLHCsWQD2/POYdVfqCcGaviN8dvc0McezxL85LqahkvsHG3zF/eHDwh/zWpz
jB3Dj3Ic9BmMoCuiD9mP0vXS+jdfpZfPHSN8hsdkpbJ6EHP/pqocllYuwE/SLGiF
y6eH25EMoQqFdKXNWHqm8+qscMPPLIshJFInLdkTw9jBt60bGVi4ahYCoBlrqsMl
WSghmHY0ENJRWVS/ynFfK2W1okeBtg8cxn2k3Xk3MDpHV1NRuskvmc2Exx+3pMy5
ayniHmA9D5RRgO23DekpXf3zo1Wspn14SBDs7L4UyRyMRrRntCcP/6Uj8cRcsItJ
yI75gZxM1s0oi6Yel37ed1yHPd//QAlsVA8A2Kx0Z+XrzQsaLCcGtRkxhJ8jzJvR
DJQNoL1rwBH0u4VeJ8WhUOt0A4i37NbFQPat828RFgcVwc7mIVeDbJMf6/ldUjBF
iw5B4ysJAxyScI1fFnEFNuEyvkXlH9ELtuV3gB0U/jtgfU8iNrw6uqB3GgKH6BBN
A/Fu/blZymz8VJ4F7yJXS9h6Dr1yAaj3nMXE7n/f38LIwMwb+iozHLPDRB5L5M/V
e/ZvWEVut4yRmBxO3rfUC9fO0Y9zwJIjhxhOwztFweWeJm3c5FENR/vjXzluURlx
dJcpLuqkVHv4c0FUiRhI8KAwQ0NMCaXL2nxM9R76FlK1b8Yf78gq2HoQNBWMHC5B
zUcGPZdYlVfn3K1fuKsC+xw8YGqSEbp1/DpJU5XJ3dut1k4cv8kKprFPsMf4SF5k
5pS5eplE8f4C0t/dob4VbfQlRechlPiYX50dmnU8yHHYJzS+9DBKOyfkSoNxmu6g
mBNpgBH6rNx8COvtvtI2WYkoHjqu/uMZaduxFK2elCzQ3riv9gEHJl07cgfvMQUp
PqJJVNtGuF8ML7hLj+mcwJgoSpc72hT6Gk4iILE5a5D7H1nZQxnUmF2UzWkBuQAg
pYaXqPTzMmyI/XI90pXU/f8FJzY0uTxVIWrg3Kid4gRtXRs4OwcIvmnoNIW4TgIi
AHqeajdCrqz1mTqSgTeTZsaYTUX6WLB5PF22KObkua2AS0rCKMv64FD9JrYtRQQX
FpZpelmFAvbHf3wJB+GMTkIifnK9jBa7N1xv2atWbIuz0OSycSFo3xvv8Al79Z62
6kxhBUX9atGbXf1qbKdaqCrBnhAmvvTMf6kph4q/x4QvAN7owD1/EHUKq0zQdXml
ejYRU7RU5ZChtfIodj2LdBWG9WLTAu3lXSXx6rB/nHvFr4XU9IKK2nX65G/AJM3c
8Y3hQK+bQCOcXimNW5cQD3beiHKq9qFvk/4gCqn2dQvoiCJsPOYkruvuP7V4ZecS
NvQro1IQG/lP2I1my02EDhaqOgA1R6VAHbyX1QL7AAifL0nNV1OX+twTJyNu923m
hz2zGEfs7mlPR6V6T8DNb7etWyJ7Qf+k7Xrrr+p2C9W+5T6GyCAyJkKdFfyl9+Gy
vKaisKyWF/cbC19Bbcchbz2D+OJ9ZZ5BWkbN1JbvALkAchF1jCigPZK2l6H2VoWt
dTxFDzzCNYtNng06ilgnrzuy6e2IJZcn/Ua+UAoSbuPj8eOszpkdyONSMFAueqYl
Xp0ZPp0fjpoXSWQsYIL5oC2TeuSucEJS+vO9eBm9SOkCZFBfNsZgq8maTBnmQ0E4
lp2ab+4IBYxpk+G7UJdxFdArtveQFGoqtbzLcL3bg6pwmcarN5EKK16jRXUhiH8z
ZiCf0lOUr17mkiKlkH/qEAUFRm5SEkxq4f01dPTfyGk2kcmVqFSLIzfmUnwruzX1
pdXTpPldEKtKBkIipGp5j7bDoLhwdbAyAWCe4VfKL9UZ5XT83TWLx2yqSOIFqxGK
ZeovQVz48eZkwdo70Ehm7O6ksacwScmPGXwaYm7Jk4BWhr+ia7TTcKDKyJxeoEy0
0ncL4bypBESlkZrZ/U8VOb/TURcQtyxF0OdafGy9hL8OdUMz+IdL9ATolSbiibyV
a5Kfpf0AyneyEidKfqQ/J4+deJObx2hHP6ntHIFfI2LQcPCwufLTVeshuLqWL6r7
2rKSWcjEJFfWkunndZb+TpK0RVRPJ24T4aY3cWS1UZr/ZX+/jcZ1p0r2FuE6nxkh
rvCbjd8aUeQzeLo4iLSVKCca0t6u8FV9fET8gn1RWbrX3LfuEjFa0Xl8VAsZCUnq
Kll1CdiY+88E0fw6GpeEr2GGQCfr2E//aWGZf9gAaVDxmopjIC1COXbKabyFgsgj
A0zFd9yBuj0EtYRc9wQLNsTDlZ+Q5JHML1TAUwaVwZBDljhqE8UJsIBujBQqBl4M
6MfxKMZG5RPMLxmCHeaDtq4PLoefpJ4xQPqfoNKPR46litDfoxgvhWGjRxX/JmQL
SualE6bJjNsoIKWrwMlbORnvB5fndpN2hSf3hwGm0OX8l9DnUdHXPwmd4lFBidzK
f1R2QV8LX6OBy1aMI1Xxsl9fk3oL7S5TGKjVZI+n4gPx2LGMwUNv8Rt/3ulRKCmQ
AWgpVAD1UtsvkY0lmw0lfxzjC2CC7LqzpDGzgl3fIi16j6r9Hr/IEQueEw3WiFEd
Ow97qIZbkl+OYX46OR0X7ysWxaFtaWvbYa0yFZDo4NIkgW/opoe7NCeP5qhAP2sy
Sa/CulalgBS885QTwcebZKwAXHcsFIzZLAKvuRNSbFXnr7bVwjLO3uvyLRMatpz2
L7wEA7ONXLC/j9fOvlP2MwB4fMOSZyzgyfjicmQFVyh/ldjbxyqO4eiWX4GJ94Tw
uMosc8hdcpZN8P6HoVb3MtLxjxJFAEp/hmuMid3bZ9L962CECaqDypZGxYIST9/s
gqT/Xr/erHV21S8Or3mzKz5qQ2EdrMHTtRRtB0t1/uXJKTgyvjUMxvqXPjjSIUue
G5oWHULeYdDLl7M5TeXZiMYoUK5EvBjIPHi+dz0SLCq1jlT6yi8P11QduA9+2qwG
vB+GOHfezJvY0jI/9hoNPlbbCuJZ0MecX+68O3rJ8svHbDRajMPPOQFsegh3VeEm
s8vvB77Dfl2zcCgrYCOqkWVq/8MRQdI23+mkqJmgcGWqFcWUuYji8oY+IhD/x8Yw
ohivWUH+I29sCictHbvMK66hz1mb3yl6m9ILKI+gnhgeuSDje6ri6vD3O284wIdM
LPfTPPZOKCaUIoIa2dgCp6JN1DuoLJs3OCvrPidF41FY1/tOoweKA/9K06DSLHFS
J94I9HuLEIGk3FjAGfhRbJnhoP2f9psD6lIr2cDFgbEsuFhymXAHBN97tbvfingk
x56Jn/w+HRc0CS3mp8vE0sAcg8+Nqycm8HTFDYYfXndAVNFfTo+o1Xl5hIcURYK5
BZQ0DhukAPYRuaHy6IHB8XWZu0UuJX7i3S0usMbLHDlM1SNyRtMKpP311T9C5ni3
hO7qeozLLZfFBUiJyZO9rucjIgEi4YMvun8S6XNcFxrrEQCJq8Nfl6cIVPrXizr/
liEaGj1PU2rfhSN0DK+F0tLFeyBKJ6+6Y6lCVXPinR9ke2f5DvK5Ag9pVrTYVKcc
iVQ45oP3Bug+BWQYnwuJECLNlcymzHdTWyKAXsuOlBHTlSBmd5VMWO4b9lTd2igm
twhnHLcKU2aI+zByqby48JBvNYsUxbmt3DegcOZwX60TF359tcLjpZlwodf39OC6
9gexvjVUAugMe6Jjx3TqWRkETqC+TrJRxHRQNYnBXkRUI5hv4rICiej9F0vHyG17
QXDyGZpwHhiKPS1oNCaVYVFmLbFhXsmo6/AmVfnXe8D1iPcM7fvKMHl/lQ18hhb/
/BfJqvyDNlGZxVGiX6C13ZSl7p43cSJs8mpAuRHrNJbA7BlW+AaT1gO9mrjvfqZg
ncZ5CyDIpe4zmB34yn52E0SH1CbIYRpVDJv34/q0g7VIIpsw/acrwOQ+MWm3O7i4
OhsomxdTSJH89qfn+9dME417rZHUlMHOxYdlH1lR0Q1D4YWz3+ifm2XsO1Y/Ckqv
cwExiJ7qu1SK4rdzvoaJktqxwYUa7AnY+Ee6Dg1cBHx3Bri9ske4wl3Io0N6LirX
20u/tb6e0j2Q1vm5yUW+Im0gr9hDxjQ8i0IUq/MLdZunhqYVbWLW+w2G5lic03CL
pKY3iSamCiYa19lwDPB4MmvLNLpXFIAspY+CEny2VcIQ4JvDKW5GaP3fJmAzpzQM
hMrnr9EEsKFD+0rH5zZaBXMR/wagVlTAfciesbo3uH+m1SED1oqR9t6oRBf6+7GR
1r5rl5kKUY3rD4QYyi9gn2PXGKGVtAPRmEVtf2Mu6kcsXkftdS0jat5P2xzEZ7hh
9Ar7VQPoS34HL1RUKKD7OTmvnagATIHo+d9s/8c7wdOj7QVZHsjYcVa8zL3DLQxp
d08WQ7WcPumo/4pu3DwghVTyI7ZSqbdZTeWxaJQtKLF8ELTytuEo+RQBiM9ri8Qk
+4VGYDhB4egnC6MlPM57DXtnxxq5D4Fg89CgzeNXPq3aPudwwTm8I4RyRixw8pnl
2XnqhQfn71n3GZRx4SEeFN799FpYeAoc2dj2rNs/FP4oGE2E6+njgtrRBhiboxXT
3bRLUOJTqasspp5QDo/Rm90ZTaHkueVpf5fz7uyketIDd6JgbetsC/+U7ZCcwF4U
q4PwOII0eazoZxsXH1AVfxKEQxDoHsh6twTL+tmLlh+lju2JjBo5/TQbQySPrsRR
JsMe6ETVT9rk/WQidhPHkKKEW6+jlP54INKr28DWcVEZS0cf3syc7SgjjbKN7xNY
zkRHrNfGMWalSuM1R7yXYi3EvLfJlMRQol6rMKFqrHtwb/DXPBSVWVFil4wOWd1g
I54ZZGynZM2Ggv0nXZtq8a4HwM2GMEZC0Cd1I9ipEfHeJ7eolFVSxp0qP9MifgFU
d6S6ejhU0gYWdvEDysKOX5uWDggumte6CUJwW3h/01EjY2ma8Nk9AA374sxOMIRf
ypFI9V036vihr1fqxpsVCFCanacSzTqMB0lIN6UyO3dYRBwvbDayvewiEcoMKorc
a9bNhzet8IglMwvVOaYqbLERVMtXIquL9YLLuBOM/bhnjVLDmAiGtp+fvk8PLNcp
4tMcmPNd/9ldWt/01USSbQkZ9N0uViGAjSbQVTubNHI/BUMSJIf1dcY8DGEZ7O0M
NVAO0VlFlw5MTkmdJvM+dqieHucf74cKQdZq9080Ljeo+v+ngRlZwrbxwE8B2Tya
2ATH//Au0Iddp2eg0vyE6UCrrgvqo96IhwxLZgdQwckyp9SNdfrkkYZLgzYhT26L
gCjCLf6s7ST5L6t+6Pb1gjtrbgd0FMlUs4PTwM2xpRgGiGOC95CqHDAWOAIKA25J
qDvSLwxtsMjxCdewg47iJp2vu1YweuIMdUYB16xF7LH5XbDWm0AHuXWmtdMH3lQ3
NSmVdPRHiDNr2tzPZOxmh1ZGyJIoHwEZAYvqXkZCmcbiHFR1VoseEOWH7qKgABt8
D3gmtQPbKIRjtZ846rJdpN/3ALMJVf+pzQgZbS4ZnBnQ9Akx25J8spqB3y1k5xLW
hTEe5TERswtGiOena9Wne91tYZSFDZz66ibSqpdYOBUC1xVykzzF9uAW787zVEUd
LsTKbd1RPKBWHFMtpsKHH8/nG75ZIw5GHAMZs5sG2E40wopASq05bbW7rJaRHeAe
Pq3/ZD8w8ux95Vwn+qcXMWhXZsVX+/g3VfhyNKJhMEj5n4kkow9epo8tHPgoUCwf
lRIlN/R+uto/eR5tRVQ4QoWxXqrZM9Q/fWOzEhU2zXW4BSIa5MU6LI2rFCgPfeNG
FxhRdlnLURebFczG+LoQ/Xg/+B7ZwZuygx4WFrcudYJSYWrKEypPQPSlJvQ7lBsI
60gPyvHO7FDm6K5Lkq29mKXSvCwwlh848+t67owU0O/OgUhbnjHE9OaZSMVI1Zde
rAwwY3b97Va8cfp7lo0lMSDL5aGmkhrmZ1+/YpZta2OCShduWLjVVwEdp2AEYpya
IOMCDnASgGIWr9vy62RxxAPUZMXGNPzs0JwUDSBAAc3PQ5Ir4UGpiaD6jVXtzZOw
n7ApvP9iYK1NsNikpICrFQ1JLgKmZGmUES2XUPHX4fcKxPWsfGLccsSR7hwM7JU9
DI8/fqWelu+eFu0DxQqeJSdvteAOFgWnnS0gfmLMT1p8hchkgfRQ1Y2cESkpw+PC
IXaXyhQ5uGVaiQCHZXfffQbXbIPI4kMEvTu1KSWFnrYLIZbT1OZqTFE0YnNgloFZ
ImbI5W/1v09rbZkr562l+GEAzpfs/kXpoZrapHYP7uraxEUpcnvLSPP+NpxfahuP
ODBqEB1RpJ/GNlSdJGlAfDJNh4e6V/++hj+qK8corhMilS7nqtllrHhX/YL1hoRM
uPOTAcWnuF8pvkm+TADEO6Ml3V/oS9SA+IA4zBwO6wq6D5wsbJCspCPg9tzymsnd
Y1PCnKjuOQwGQcpSB4svM2NduSL8LPgXwqlKAwJMkAj+NPTF13LvthceoKqdZCOd
QHsXtwWFJVvbq0LDRvq7DfyX60BtU7EeUXCCEw/HKzEAo0w4ptKBll2VIAJ0Q7ne
B4uG6+cwH9WJLAplEt2OuAzWl9XXNLNgQxSHzq0dvMkWVIV8uIAdlJzc3RE1KEBH
nlPevvdD/Mf01svOdTm8Vxf0KnH7OSFhRm9+iDfC4NfOgJQtRbmnwCcyxFPly3pL
6+aSory9ib/Mpo79dFEIkcTIFkc0hML3EsQwm5D5jLaLnEIWG4nfGMlLQVW95ySm
vqFaAWShCNVK65o7Zt6JUbhbYpdMle8lWr1WPJBFJh0vleZ9oOCOirNrGpQC7gN8
uDH8CanFNPxLdKh1gE/Ivvm1+Z0M/WxuLN6cAdavKMQua5G285d25VwyE1UDGYXN
JFrmeBneKnANTj++wSg8HDAY/ThSw61HU0A42X1gFLQCBed8H2tJxBPDFoAXzS76
4WEXbCcHG+Ba/fRqDHbLlixltdXEkSP8QGZEgThppqn0hLnfdT6AjKKgZzfCY/KS
V3SOCKti2MhP0reJ+NEa9kaZSABPCPUEe+URU9BMlPr8Eu2sh1TyZACMAv+cOeED
U+OWNjjw2gBpLy39NkZuLKXyZrjkGP1s7hp0aQ2iEYaWV/VgfgJmoY+AOoGtd0E0
CZCILrkQuE5DPI/CsZPRwA4qlEJY18V3ZKiybGmTaza/bAtylUB9FjnTHCnqsDvt
wh78I5VPWq1r+43THPEYj5MbfaexsqufvobQjkTKbucE+pQlfNgxuPI+FHTURyw9
/lXy+heS+ZKMqbj4a4BbCB3ACc1OVTKuHCy1jbaSenX3pQ7gsH2RBvrVVOjkR2Ue
avK7JOjvaoNg4p5okf4+mxd34+rmGNc4cUdp9+qCkj6jyzO2bEoMp2No0AiQENkc
Cbij+HDwQ6i5V2EPQDZdyY9KUyKXp9099rXWbDweUh0g2MqbUftMNPO+fAjidSrx
/bBgTmVLXGMjz2/ScQfhNRqOqKRu3PAiMnMjDu/Sv/3TuPtdy2VYRqR10SZFSKCz
LvSOUqrtZs7s58/FjVXbf+wGhwCrOW8bcYvZ1fq83ephq3qcvtIwIVGuhB8uviJ1
Gvr5k94EvqdGJ9pU5lUcBXoWdkG3UL3EK8GKkV0rMax1LZGFp1Csg10+xwxv+wvU
ojcZ++NQKYYLiSHFCTvhwGbXJhSOzhdJMCxONop2+2ezH3QKOGCA2F5yaJLiuY5u
sXjJhj+0c87AMj2we2RoDt2O1bWGcFWtaVD+2zjJgedB9+i+ADnW40OGBgnMkKms
0+a8scRFg1WU3yk26CQOTPBffT4Od5hKcXA+Ofs1mJ6/+M8iCQAVe8Y1MIqtslsH
6CjeSVFuHMIQGKUwizyq3jnOBEdRbpv12WeAwKdqz/LUICBMNNgMUTQdX2Dh/RFc
4rTwqQH+wboZy8yHjS6ngjMU+VnpubB7TVPGg0CGlivJA9VXP4tEAhxQaOmFdjiK
0u3lPkEELu0ixxh12AYUKmITl8g1L/tUCt6sSkM8CTrFogWZL+sxv38uCq0y3x7f
5CLcWk9ldTcV5kJKEE/n+q4Gingkk/H0+SP/pQRNl1upl2HsREF6H7I14odPELl0
ZaP0w68AiWNZ6evGjRC3irWX2HLNbjfvDtAn10K9ZnV7Mf00VucePrNWfJgP4B45
fAOyo6UVH4eBPcaQ7dXnGCqoIFcGiQ6pmjWEgO7KCxY8XurJs7HTFZuKgfOCRTQl
wXM/7sq364gJruIzVbEq235YHO6MCu1sCsJsoGNLDIATX8TXb/2hYwEmAymyG/66
+g5Q5o4C8AZtwiZZStnMf8xCcWx0tl8SQbbxZKoRdyL376ha89zKjU+tt93VKlgZ
i+hUap2meLGk8nf51ua+4hL9DF0aY654+Rrk1gAJd5Ca+YgPa7Pz8l3JJlG1bNGi
GB6Vl1goqFy/4I46BhAQspPPpVRdLc6wmfO61preJF9stZ02KT3HMcx7jf4HL4Ku
fh6jXCwblLj2l3sOTgAsm/WLC7SCSqz1VLY9rr5Te8VWhUR8tKZc9+IaqM8mjo7l
w10wVbaAsYfxtnHTKUWFpaoguRE/LfTjqknb5Ck/h0dfalb4eGK/CoE1O/RxeUic
GA2Hi+7WsuWypAPVGooCnZA8EawWcxDsVyVoOUrCHRv0FhnB+Td+Z9nTA+VgxiO6
W82US7w6wxtn0ruRpjqW2EnoC5PNqMmSWr6dHJF4KxnnVj01nxwXm5o1AbMYLX5t
Rb1OAEongMs7PwpSLMkrLpBf4xm/tkcpYRFnRaKT+YlW71TMsYu83k8ZwB0XwCeb
3OIeznIJ9dpbs/XX1X09040yt47y81aKLur0oPQI5djTYYB/y2sa3SynhJCD1IzV
nHCLqipLa22XpsH7t6fIDUJEJkinU/QDEmoX5bdBtaxeqfmNRCtgoR8mWsti1pNz
jRjbaTYzwCiKju5ADOhWf+lyYFlFaiQxcdd3wvz6qgaF5YQf56lIC5t+rlF9cZOV
z1wHKO965M+0RnD5oCdQWy+xZZxcI7CUghgbyczq4Hq+OJcG5r5NVvtpvDJr8nAj
A3s5R8BDmYwt/BAvhZKAY8jkzemKT8NYAvW01TDFvWRqdfSqfEo31XWjtds+PHw8
q1oHWPCTJrvSItjsGDA4VIiDPouLUPbofJtuYFuBs7P64MwJoD5FgV6CiWQm6rW0
wI5zf7CN3bFQvTyP5sFpaokLPQ6oZC5TDJF1Pz21tXhCKc2HcDuLlj4tOgJEbTDZ
wrJdAnJR/dlCzWBW8z1eueJnc9QFgG4mmakz6SwEZY+AiNKFhI6XLNbT7tyUACHc
68fOL8LwNigAxXxQ0JOss7jPaFa+7qJnhd3IP6l+kjXx/gDX+7eJHJBaXTWcn1Qm
3NvUlZthWCpePthU6/unsuGrbi6+28u/bn/x0GJe2nMKvYHhTV5QS/KLrt/akWlP
WrX62AWLIsFD5AVbZwnEjCNCLLvlIzf0ekY4phu3p8m9rcDAhA3nvNfxlbDw9VM9
MFKkUzTyH/8CQf6HavNHbEmMin1BFpWKvUcm2+RD89qbG0PbudF122NOjiovFdMx
fULtQHSkZnsLKyQ2iVC0AeX7cT+boP8DKQeai4Axom+6qLTwLQRPTmRHu0N8TuHh
Q7c67MSwQiHxPUKwcKERozSATY/hwliUlZYCFacIB7P5SwPB+0fIzswKME876tPh
C+rOzyNJ7xbaPv//JOOwKztdxKZXDUDrwOQSTLtroHt+EZ5xFGCHf+W8WeuO/y60
ZSImo34pqE4KfO8/vY8iwITAnszp0diSYlWUdIkH9XDZ/44Vwz/UY6ljbnPfuT8C
xMP5fYM5GKYz8B6eO76IGnHFFs9vKnMNIFenROFDLQOZm7pu3LKF8QhL2irftJvU
+Qoa9f1dGz3EhU1NW17+Q7YGwiJmlmmc+lryfKXK4k44hzPPlOmuhfso39Tmpcg4
oBksGUGssfhiNz8XxuyoJVkojC6QJxrF0y+9Yi7ipoILQVPNpcocqoZyyB+G3UP1
xrrX8g30YIYLIL/fz8tc7+4TL1iYVl+XeKsC6EUoEd8rOJ24vR3f2DSW+Ph00M6A
llgLVwJgdEHcdl1IHQd0SppRTV8nBxKHiY5qy6hymR7FtecZJebMG2rEJJ0VXu6c
fbycqvgUwGfCyIQJ8s/S5Yf5fdA+SNwi/1nao69Jwkq+gxMIr0N6D94ZlENnc/Af
VRcryuzvflMDX+egCvefXxtEyO9/AWfXxj+oUxt9zlgJ2IxtmPe0mzaLuhDgstTx
LilDl/O3wZY0qB+uTG/sjicQGvD73jLIv1bp5FbWna8yL3m3zaTYyLUWEddJRx3u
rl8yu+emYceHK6DTh7Sl6LLUz7t14iI/Qw66cISYOTrb6MReKTWTKnC+INRKp3lP
vuRqJMzWLOGnaWe2AYbogIEGbZDASMSbMgkzdSVjpFAv50EoT1h5SONcV/xpPRYt
11UiMh7PhTNP7AlThHUl7dAoVoWRVuNekW+imFoL11FiljR+2kxDgPTh2lIqPUYu
LyK31tS3/XvYdlCzn4oO5x4KSMersGNj2O67kEq5cQNo0fSPbwn8avuss22ujdk2
PAlR7lT+CbGRbH8SqkSP7n7DYVw7eCF90GQFyqwioN6zsKibYH9BitSZ51tRE6p/
SxKB1+qmdTU0E4oaUony2+s3KAxkNMS0rJqMd+56lPE3L2rSgPB5WEPfxX2rmN5+
fUrCaXuTLGLLvN4m+85QpdFvEchI8eDz7S0YXL9w2f+yDraV0/wZVtwAKuuAfzm/
VQ2XvmFb9btbiVBGcXB3soCOXy9nQKL08GpaGGRNaqz95vX9U7E2CYqslof6Tne8
07isvn3bNZt6WnnTmytMKFx+UdW89+rfujc8PbHN6IYu4ogja2PKFADlVPmFKgFC
TGoV7sC/HgDCn5NsDLs38ua6QcAwoxmloIEs/lcMWTHSNij3g2FXOu2jBAdr2/Yo
t2B+vMxn0RJAvsaTqxJxhyWNyh/8BfTxNMtsf7kZsGQ+lZRFZ0Xag3jAA7+fN5rM
axj8MrwPoCqcYojkoGXkRfS5JuUV7+ivDqd+GOSiQyl/1ll0DrESEMNWUabUf739
4Uq/hq3BdGzwWOwhHirsL0Tq7fykd/J1q26tjOBSW/kxnnykAONz4ofSI4mnB3Kr
IGzWw84bRKZJrfclFBrmLcQRA1hxuXbRcyf0Z88rQmTKFSybJMPqmqJAmonSg1CA
HC6BFmF/MeFHsEF2TdzM2nidhMQAjawcXCzV+9EaNrfhi8P66Y6QwUmPsoo+pGGh
wTZgqDWjudPYKmtpcNttOPX+wsO10HwG5ESBxwplJJFbLbG4pUTXxtwOYOFvSeWt
wzRo1/M3R5TZ4EBWu/p1W/gkW9v+TAFSPxmLeYtSDaKhb1LPIrtsAg+CwXpIjtUb
YWQt1JrlSpZuimiBAs3EK3G+rgxoSh6CHLNZnbYFGXcrpjI9h1EYIExch0r2ifUf
/pnPJPcYgwmRMPfdjaBNvI1uKQVQqWAi2Q0V0ITAKgxAI/HqLO1/oIcfqwfUsmFe
ThxniCnFUrYhZToZF+sLE3S2u68OffgXHOls1EC6AgH39iS1XZT3NsGlVaZJlw9r
fdXnLOE66FuLNMGNw5jxwSdVDS0p2g8eXITboCHc+U2sZU0qCID3wpVvs1ohAEo5
i/Zy5rjHRnpVwAQNKrFG7eWQsdiAc6GN7jrxpWdjrPg9SiKRH+8plj29fTac6+Zm
III5rL1nrEMSTgHfdgSmFgj5s+skpBxBnqcaZpaUiYUJy6/nW91inhCM+MdqmsQF
H092K6ckBSYT1Zgg8WrIEIT4o89rHUKezLWYAxIOq/vstuJqs//gI4XXtSBqDe1H
hfxo64ieq8QK83+yWH4bo8wK3dNzcqVSn2i46YKbO5C9vjBuuXTYSewYwReyWE7c
PTP7uUnRzyXD4y2+MaIS55zwMTIZgLjtmgyudElqr3iz5kFHya8RMkGpu2gdxFg0
FwRYoIoWtiGJB1NU65Cz7TLYBV3+SuAIDRKBu45JsLtmlT1vkDzE8cI+CJtQ6Fx0
Sf+bY1+/DQV2qK/iPDpyQeza2m0LICzwe/1kgIBAoNds10pSzD6FRTk1Xo4vC3VC
T9/A7At3M6b9fCL7HM1UGDGwNBPUZG3Aav8y/Q5PWa3ZBDkPgZwltOFbogWECCzq
m9O0nzAu3dSzQsVWZPEipa6INNV+a9Y8/MqBaEny/HYxF9bhDWA7n8gK4V3T+nq7
Ad4XvX6WiA3v906iEya+/4tCKJGDbUH82uz/LXXuVuR0DQUwhBP1IvdrZmd8Jt9D
ZSdjDq00CCaQloW/LS7RVP/fJSq9G/RW34hkwgckm4IlkgAZ9+i5vT9EtUz9Q8NT
y0XM0OaYEmYNKS5hsTk6NzG9rd3dCn4BVyXxwINY2Q/5zWnADAlrISE8YyYOM0qi
l7yO+ueF4xDHrR5xb/QRoeB0AcYYXpAuDnVXFFHSg+mHZQBRAT/EbL3624jFbL2K
d0b4LOrbXLuYrOLIga9QSAP00yvHHGJUBK+LL6tWtI5cCXjAD9nLg2Zwa/YXJWUV
kV0QcqhRWPHk196gu2PhhLQyC8Od0TwhlpmN+NlqBfYgv4hqoVa09ywvyswVurz/
4OHqBF0Ix0j7kwdK9Ygs130FFyk7b8GcGj5Laa3l4c3K9nVnnD2LKExyDWEb44ti
bjERXsxxQgMED3EhxP3YS3FRlZk7WgjnKhGD712FQLD1xPn8S+uXVElw1jZrNme1
tOGl8sAoz3akMKbErKLtO6TNrWdE/Xu49gsFhbLumwSJlDP9tymP6s1lzVvVvrGH
ZSV73fcL5l9W88UYHrxv2sBOBBiW115+Pb76WkzOhPQVYlp9lJ814n8fUvPzOnWs
TR++YICYqsbJKekbnHH+wIAcd5auV7QdRLHD2sii4wpoNms7lVTH3gwGR54F7uST
V26moLV7YAtnTX8szoUZPfvZf/veZbOH6h7H+I+MbhHoKc+BiEvinAbiYXQyxLwK
cK52JhOH117TwuzJecrg2PwAEaRd3X+7N4Wet0clS5ta4KS+j2aiPFmg2UAOoexC
Nbv/VvEO4hA3ZHpCdA/TPtbcAfFa6boB4UGzTXUfdSdWD5/rRx1mPts7HLqm1Bcz
QWI7OFFcn+Bcr8vcCgKRary58BXNYllBgxI8sW/H4SIrnHQguPtvp7n83nFSTZVb
lYVfRB0t3vhY6uikbBbWhlftE+P4weyW2Y1YBfKaNmjDajgrb/mW0E4M4xi5YqXK
wCSWbBqMGyNaQ6er2YJByy8rDQ8bAMW++IpzbJokxd0Xuy7ZERUEQgi3e5coJm0l
0QVshNP4zkMaTE+2bii0kDCWks+5O4AJe2U3gG+vR90XbqU8+ETp84pMHvAMpVfZ
VchMCWyEyU4gAni6RayT7A1BoBzp0nRGLfqSs9YLCL/4rTJLHz/dJZfuty/0ZXGC
TxCnTZGNzAYv7yhTHadQdTRpGWCBsO8tFjmH7l+70jqXVhVHBs6TzlY87q2LmB54
X3Igys9URyLIiFi20IKp6Vb+JvBCiHO5EnBs5Iv2TddTGOaaUjrtMSkUx+KcR6iy
3lFr93luoqfyShyk8NarvwEpNZtXMWXYA//uND+edMnVIfWuWic8JXcJGbOMag8c
OBrjGdYZlfL7xV1rBNlki3M6Ei7LVPjlOQDn5mH/iFJw7Ir2//BW01V7se1sBdfM
qhMJsdJpB6tPh152F4ZKDH6JfC4wTauQZ4nzEsnjBkojOkQvhz3S41sf7QzT2hGD
fkRS/WOCjL23mfJAJPoiXPTk5zw9vzKg/TW7sMCRt1v9ta5sBDH4y4op+C1TcL7O
NDsz9ReDzUGOivGr3emxikhjxi3/t2EXymvMHVlEcfxATSlrJtrIS2qhQVyIQcmI
7w3vqc1y3MLY4ktQMNXGzJOhFyJHivuqRIDgGqSuGIH6U/nMsATD/5f51vXRFlQD
ixB3X77NKm92i5fkc7jCM5M0nTTUve8lhkoUAB14Z1IIRG3Df+Ns4I8lqQYUWpEi
OEPXfyCFnFvnkzhwJpTzjXTYSV41meia5BxDvtkwLuDMvQNd5ZQej7HdIMJxlH8B
XVrf8rxg1WaA5NGb/gQ7vRQmkjIlZhsA5BohyhyC14RUx69/JFT7cUKn4mUdB4nv
+JriHAixZYh/p16V6CmGNSbG1txlJRRAyxAfAW5+sWPt9kl2C/zK+MJAbYOvH1xq
3clyWx7hxZsISd88k9+KUTQ1RpbWs54ccKxb4txPN8pJlucsn6KyEkk5ou4aw8Id
7UPX+IP4mh8b1WCz59igFaSktaZnANMziXGaGR51phJnDBE7fqjR/PHwnT8h8V9T
N1emhO2039JL6jhT5vb+Odr2f3SQdSFd70GzDolyxQLbZBWyxSB1y1ePN2th/SRQ
GwcJBWn1jDa5ZpWGC0vwppGkuNdSRzdkpV8fpq58CtoiaV8whjVz86gQgWYMxAxP
pglVoJexUAtGnouvz/ikApYeAXoKtC1I4ErvA21AYASveVG6c29AfOzRN+o7aYvv
sn3c5vAit1qAI4blefjTguiaTNBK/QytmztXZUlBNSM7ZcmG6QKxkbhpeAXYWQOE
/HLMB0t3iyapxsYEDMQ0wziboHGuYxTaJT45vH/WNOavUY2J+Y4sYDuZDOabMRQV
NCkHFCWGPNaxW+YD6o89hlJ12hUJc8mV3qIB13kAq9tcwEZoF9NQ5/T0mPYfaJgg
QB9717xhcQI1PN7MEhnG5hLXBM+Y+IvRFwI0yO+sG2b/0iaUuc6pFQX4nv9QNBSl
GeqvkzrlfDKBDI3KNmWNEJAv21OJNrfNc0mjE3LCJ4CXUyXPU0HYnhj55B++bNKo
wxbhCQYiG9H6ZsM3vEc2FBrMiPaEQIl6+mlqULdOhb4Z/iGQv9Yed1P47SX3sfgg
mQPtTUyZjip8GS7mG3Xhu7+OP5F0kDy+sb5vmm9d2CSZa4vF1dMZLjeo8aWIFgqW
0o1LblzJfDYoryi5jjq30Z3FS/iDUR1oLLPKMaGImWuXdChBHaCpZeoWBPgzVOGW
zow/QOZhEAKHA9ZnNPUYZWVBJP4jZb5+dPuCKol2wCSKFfsOR/Rxkk/yHht/df1f
wxHFslgZxhyFZG8FREsw1Ak8ejU4N/wiWbEigeYTHAr4Z5/S8Dha4QsxwCakhiT+
qCjrTNJ0NpI6DaRdtoeRCsU0enrlpnc6eH1lO78CIGP9MciabwaPyzOCveczFOwR
OZ+E9yrBcSsj/5KKk5zQWl5K2JTprxndITmsTCIJbr6tFBFTHKO4cgHv7kykcGyR
ksukYV/Td9mIrdzvUlrqUnjdPJrr/+KJ9GpKplO8G5WRNMyhNLW8MnZtZBO3k6b4
YweCxDgblzU7rSNLOTvDxGUU8CwLQV6Le6CEVE7ceW6QEuoUiB5e4jhCNTUG+KFm
Ymgb80bQQ0ZbZNoAUDtMLiMC+YfUJPik1aXe8n2HX64SI0MKri6dE3SzL6XUI2TN
W3As5IX7qybuEnll0Ub7W/G9W5zkI/Fo42ulA1ifd72W6SSZyhQXeHJUhyqRErv7
O1nxMfltrIYYLDkEUDFtAfWUYMpOVsV9s4hnZjEB6QsjAIn8HFmLHIKQRgoGxZ1r
w2uyKXSKsMq8DQ3jUHY45biszMhEdo3mt6R8cf/GZRKZhzrV6BqbShuzTVWAGSLm
FGBZXiw59MmDtijuFM0H/iKdtn+6wKxo2lomrCD+fl2taVHH7tq6QJeor+Ismj3W
odGXeQ7H0r7xVXOEkC6d48zSAZaeVLcjGq/XK0LVqvynOto9rLQpsb3zmGirPSNQ
ISIHYO+Emfp91khJFIzSK4BDGJkfWAr1OVbk26PjSHeccLgwC1vumK9GPgxENci3
OwGTJLP837Ey6wGzR2m42rQSkEPktFYJCboemnIL7JJlfSWBkeK/19csl1cKUQcs
oM6LE4ialBb67LRryPsDHNGI/Cr94vswkQrOLwbYfgm0pWxKL+Du33EbrJVZ9L36
iv+0Uuy4fy1Q2zYwlk8k9G2WD4Rh0kgmk3qasvi3e9pXU8LGSb6wHLJUaYpgfytV
CLrS46Wm9Tpr4Y+mdR+8wu24aZwZYMWlFY63XP8FKpEJTRPk2mAtXdEUVme2VUap
dJXmAegQ/m9FAHHw6VbUNUccWH0NiABHYXE14Ps6gil+VswZdbeSZBIPHeq187kF
HV2egdziAFaSaanQ2oDUuhYlbx/MOtn1WQDnL7iHkHYIUjL1a7zr26nw2r9TPgv3
gyASznPh0I7FQakYmIGlrlskalQfxyenrK+aLjpOdfMXb2uSn20gqI7DaREJ6T3B
2zV22TcxBQ92UeFoIvpdadJgqmczGBsE78JAaZQf70wUiehRqxzCmGpMA+cIosPj
SjYgHDaQz/+9MjU+C/UkWRjVZ8UEq1Jd1qV0EXnm3m10mm80fFqnbj89BVTjkc/3
MEcBXZM2AgLSkVYEV0BvNjSJR5PdktMSJvClM2QHdkDDwyppxtfl8fpbYsNbPUMx
zk+OeqLo2y8ceZjs3iYOGTBIDdDTnDAbGQiXdFyrmy8zjfS77RtlKw6dETuOV97k
2iQJKa3jH1YnCOKG2L0dHN+uA1Iv7OheSt3K900lCBQOmvgf95FdwtX7n/xIvE8q
xkX9zTJFh5O+QXDXvtcfYLx9g1t4ZBuW7cGCbZ6gsIHG9ZvkY8FOb9ghkofutLbN
HIAYXdB+W6UY9o6G1yf1qV7wrRh51yNXWeJIgZwLwRbZJ+zYvuozMDHL5IL/nN+F
CuqbYXj8yuTg97oPeM381J8PQMmkb9yDrhpniJpqWa+v/U1DBobtYULsvwh+IJKg
8rqvqMg+GHS+5G1gLY4Qx/6hRuSwukmNW5V74ilEOQ33Yx/7IrVl6oqAvG+pVfer
ecpNiGrHkUTyTg4PDvR0lBldzBVkhfKymUSY0AfVNBoFaH1R0TesM3L0azGUkARM
XsKbq5f42srcwX8bzaBg964bdKmlnxrVBWAq6+fm50TiPGIjRAQuKOei1k2hYE2J
x0pJvOU263WARBT0ScqbAwoytyK2qF2GLyE01zKKuymnyHjMw/MHkFUQgALBQWm9
eNOKLeuZlpj/hY67BXOfgtQm+u3FcaKXAn37HVdIu3HhBfjjDGj+rWB+mBAjlgZM
neXSeSr/zsg4RuGLVjhaeZlElvPzF0NmjEmsMSZpPkIrZkdKgUk8jEttMt9yc6U/
q5DXp5bcxbtPhsGQduur92L1dm68t6mROLV+YQBWJXvTwwHG+mbOoA6hPdu8Bv1l
OBMgAlldxdOH+5YBdQ4mD5kiqldjJAuJ3WH/GsDlC37mvfo7l7rFKvL5HmpBy00M
NtW+BG4qdLGkC0Y6ONaip3APp4zpA+hpq3VHxDIcvvPtl5vLpjDRpEN4jlnwhNm4
6Iu41w2glCS1OgnHwjZWAC/+cSLdhOznHQqXjWqCdzcJmmqjStAkFHBDRG78wlZ/
yXA4BJc7pCEQtBkVrOvW21Nd3tEv4fJ0+hWYb+IlEvOAzrltUpVlfggBGE1nm5f8
MkU7qL0VZXNZs99MvtNdBRy8XebqfZChOqX6wGa/Euljf4QoupC/6HoUme7L5ppg
qHIJ+IFvNJxsY9x3XMKaELq8/Zx8imE9GEHqFUP39OETmgxQBso/Zrrk//bYGjrl
`pragma protect end_protected

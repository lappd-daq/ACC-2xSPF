// Copyright (C) 2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std
// ALTERA_TIMESTAMP:Thu Sep 13 06:37:01 PDT 2018
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
FPLotb1DA/YB99EQifq1KTwLDdoiutbtjWk4J2qkCdKEx4o/mIb/OC9q+gIyL15k
Kobe2vFX/g7Wkauoi2dAdW65+e6Hqa3asXFkDd5t6SOS+++G9UE1wkmXlKqCH4p0
WHnjCZ5UnQ8jgaDh3Qcywg4BMACDD8danb/mB+o0UTY=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 7920)
EJZVNBrO1f9YHKunlZEvz5h1C5idu8kiGhwsVfAIE1TKXF1gcXAzx1NFgCiBrm/X
3MHjsT5w1TWnkPZzZ9GD8XnPPUc19hKvgdXYE124DF15QBjT56n9k0m/kH+6tQM6
kfKOTtRZJeLcDXqPJqjMf6UicBMhhnHnQzonP5o7RQJ+nG281LQD5P/SGsLQtYD8
GfvYCaC3QsWqOR/8Dx7BzolIqZ21Oy5LKn3RVJfL1YpOwa3sKd7ThHD1QeQ83dbP
p/wU3P3It8ztkAjQQTClMGocYDUDfrXBTiz2QvBCes/tBCnUDouwiFK+tU8T3EM4
/46Ji7eprUObqlFDBqD+/tAgP32hrfqYHI8TskkuMTf7EifQpMHrMCaA26T8S3VG
nZ1CgknLRdp4vHT/PpOef/lO/N3lAHK1A4ADBqt7hsFOUI97nBLn650+uv9cxDBr
hfMQnX0SxnAO4ncICEwuPvc+r02b4xCxefCultGLEbCZzr9Dgha/cuGgMz+20qky
4NGBD02AOP/7yQwVGpmAwmAcId/+yl0nJtd9JieaXV9cqegCYf1w1JAxUh1YICKL
Nxi9S3C6AUAhnAvwKdstidYQ5DjjhkuFN55CNwNbs4I7a3SFCpCI+GRlF8yt8qMy
Fgf2UFl+05+fa05klXIFUtzo4+eM87eHnMmKzpjRWZvPzh0rwRp1PXMwWc9AGaOu
Ap8mW0ad2YuaaAktpYwuioDBPABS/AKx11Hz+IN4zDG6C7q/AQmntO4bHQPdT5Yd
kXNTsAbDVfHpS1H1bbFWxk4vnamuG61of7bqsrXZtq4g8yS8sRjdlQyLTB+kXxj4
5qsbgUrIuc8yiudNEEcTKmRpEiMutBa/3ha32y1oJskrdcs6arn4E0BGQMI/5iwy
Bu/yHSfOnvTJ38nSFFw0lbj3fMwop91bfgmrgcC0zz/t56xvT0kNFSZcSKreRvfX
x6KerT547K0DOTsgT+iKyF+Od8k+QLapGkdUtDBozdrMbY1s/EvuK7YLfaVEx034
4yk97aJEiYQgW8t8aqVjKNGcfbiWegMvFQEAT4rcMtiCTfZHxYiICtW6kd3oNlfn
7HTvB+Wnv2kly2UCcH0e441hnrluVpwkC2x5R43CMGlLvLZNhFz3juTtw1IlNDum
OJb5nydiiBV4iQpdi7Fbnv+bjaGtm6eIqFVfScPVpv+Of34c2GXrXTEAQUSJy6iJ
tvGRCVu3CaLAROGcolH33m2aGPhgFr91qklsrUXknXqexXlhWpH+xsioUvmorDSC
rHk3RUdm05RULZL8AdruBXj1t1SPFmZOYtoYdtj6pDCR85BgXJM64kMTP6Xn9PFt
OFmCMp03RMaWkxC06GlHWuGUZ8+bkK2ND2Ogd1LLzQr5/29KRVtzL/5c1+ukdvL6
CGTc4Bcc7EuJTOR9vZYV7+wMxqtizNEolJ1CxLa4mgiNxoYLRtrU+H4sllAYT8Kr
N4LydF9B6W+XdZ6Gz5Bzwkuq649/un3Bn/sEkmvazL1UcDkJc0v0i+juu9+9c5zw
WYjdY288bsjP42wUguv9NHeH6mPgWGLmd0gjQNv6gL0uasI33D6p3+QJiakQxA0X
HNFdoimvP3B96sDWmsLHk+dHWJpq8YLmiTvEPVvZ6mLbozQ0Gk9qOTqdHacQ385r
mCA2MtGhF1PzAr3bE71QDleDDGhnp0yZGNtxGMUxnEG+H2F+M/zQRFcJwJaQVaJe
fNy/XhOzyCPK2un6joXPK8WOS3QNA5SGif4vKcuxVRnxr9eh/w7KL7QGpEgHPeuO
zQsyC3bK1x77Ikbth6unft2c5S5f1rNTomQHIpB3PfzdD4nEHaOEdTonCEb8f3mQ
EVmvTfN83j/mddOJl0zlbaBnBrfZycI+BTG97ZLpI81g4qHMSVY3wz/DP+KaTGxl
5qthRiXGTA6dgdK203yvVMpTLAXa5qS1yJ9ISyImywK6rjYByjVe0JKHmpUossbg
XxWPZqesVW/HdKZvcJyyZ3EoJgwcCBUYcKosutKci4gHI4YaRfBfaiRn5OiTe6bb
nrD4/Bp3F2ZxVOUqN+WR06NPvvOWkF80t7pbMQ9CH8EtxGNq1++8epjnsKmJYg2p
nOAUAAgOETyXmneYlqk2cKWaPqR9ihi5XhAa4sLVKRpzZHjtyyrw8PB2Vv8H5yPP
NzwVuYH2JlnCJW8+uUc9+fuHpz6SYomJMmOC500mQvWvdEdNqrcxreYIAWtgo9VR
/4fJOAXigRmYbvJjlsiKbMpntZXgZZv6L0WcEADj6H4EUmHUBe0GlR4Z2DasUceS
iLUGrQgh90AEEiSmQcfAOmNz4bUar0Fa0dTIQlXTepA2OcJ4n5NrKpqDFqjTX9Eg
ATiv01bQ3rV8dj3ktVYDVZJcKEytPJG0Nyt2QUAFlbRBiIS/9pFwRhHyPz+2v0Kc
T2c/k4OGd/lCTQGOwktNYw8fQ0hsu8hmCkfQNKzEaJGzxM64gWgnh4GzklOXherN
oR1rlf7ETNuhaHfG8R6UCkktbfnQSsBXzxgeC6rEHMihLMadM4h/NQeP3pVRSreg
N3dYjQKPFs27fihcb4Q0Mb2U4qv4Ro98541Mo2PZeO0+/ShBGd3i8LFk5JfsZd3G
QGVmSIIhAIUux47WXWleVtXWBH6eMiHNcXkLFjDQxKQQ28qdUemtDift/nvgupgQ
jVzk+DIecgpXHmTEA8mP0D3GVkPoGkgX2AT1tgXhc+jW/BuWmgMOOx04F/gM/Pg2
V7DNTyBRO6RwlSkOz4cm+1STm80FzVVjLE9R+mKduWU4r6SfppooujUpALqo5O+K
o/g40qDD2wsnyBbhu5DvJ0bYK8BFbjVNmJ+7RFTAvkBrg6yqNO48pz0aQ4ci4Uvj
Mdnu9inKX/5oZ8g0tpb0WHBbJYOwGK29c7yBPB3BXnbDeZrcFVhyOvCHD9hHJuDG
6sTBA3RX/KC3dX6hS8h0862klYewQ41RcfRSvMuNq47JqE9U1CjjDtDzLcEAKEMK
t2maKHnGD2xGF9eRCxgAqZOUXhmz8NEhof2XengaQBX8v1+dBE+cX/OcTyJL6IIQ
Rmx9Zzr0mPuR5CgbrKidHyvBupjuHAh1fBu65N1lrHJQaCBrny50z7h1pj9E3+bW
M+1GPWjQX/YZw77/xIQE8MscIrky3r/eCkoR7XRCU/KfAvJoAbw/hYC+4KICKDYT
PWkxG1zI0w2z7KU8ISG7h5Huv4CMMeJ9udr/Mjau3Gi4DxO5W1CGqV+9cmb+6agc
Gr1iAuhkjQ4i64SVJqcR6ZbbVmL+4q3BAc8OuXW3Cz7Fx7EFrNV80OnA3Txco7d1
AFTF5e7lpeOIX7MeJ+jv20U72wB8Ct2e13+6FO9UaLnk5eUTyBDh0M2ZjYdi4ocj
lw0e0Y40FZX2qcqp7Md4y5ZQVMjSx2Wm0op9wPoUqCz5YsSAZTjVAunCa6XPq/A1
GzclXU5Nc+fNyb6z2UAgY27nVkpwGzdi+j8wFs9mxPNwPvk4bbbATU7OURVkk+iw
U82EwF3ba+DR9DFIExjiIsZEjWK/CpNA5hHX4nahvDE+6C2GEJI+o395FXQ+Lym+
WI5NDsfP8a0q7uOSDPcYgdIaWWuQZ/GJJJ/djAvrZ7S39ivl9YYRJq9Gh4waajgS
G/FKqtRO9aFObX2uTiuwFU+cz+6L5nUTs+8OJiGrWSYxH3Oumlj86xiEsIWXGZOC
1UqXvZ7gNdHsZdk5bih1RFywmbx/vUSRsqAe0/aqka+Z1PEsJpKIsvVlHYfmhg4u
yMtY0XBwdKqtHflyq7e6UnZ/Kqwv3Fzg2wgaxWYu4xmeAKjiEYt1vjKHTlL5alaX
VIsluZPmURT93aGfz/+wpYwHWrPjF5DSXdEm+o0R5OlTsjbTR7wn/LktrO+KibMN
i9TnQ/pWvDhp/aE5KgMnvBUf0nUeAdgi3tBQe3Qs1xSMpx/AvFPUFFsRC78Zr5Y9
obiiy/bR2KgCTFg5bPQPDXlBPPT0dB3cQcyRkr+BZr+YR1BW1isr9/sHeb6oSDMt
bCGGZkuP+G/cDOfzK5tYMZRjcW1TxqHeOBe0QZGBoDvklRKwC6NxD9cdri9Db3C8
vlGwmIafmEC8i0qlAqduHGtxZ5Sst7C97EUA414jSUB5sPm8Urs9m6MtrM1Mc+YE
eUqBJ2NZYnOczxvou7PoT9ANLdSxFOoFW3/NFu0VKEvn8oD7N1OWNzzDRF6FYaPN
woS/WaSYbPmFpanRT/4ts0dQnUFbBMpRqVeL9lHFPamQrrP/H2wc3YpgLuJ+ZYr/
CjlNHa8uC5YfntnfKBzfHfg/vm8O1cOf9s6U7ZHM9XccCWfxV+LZ8gKiPkr5n1rB
6jkc0fMC+4ch5aqgDRe0nTaFk59jlb2n34plfSATF7GXQByAhqFkXw6IgskVSIvw
bq5fhoIYRIOm7e/s0vrKu8CZVkJ5Iao4OsxT861Yt4uXKtqBeSO47FcmNEP4JW0e
0rm5sPwYnDfZMqb5IeXr6RvxGgxJeyhEO+KVGhMmlJF2PZR07YeJBMdzxYOt9YKf
8NPAAeTdFut3YdghM4mD0imdRrpmNgVrDJkXwkAy5tcaf9jJx1aQjqYxpHQr1X57
16PcoPwbXq23iGWT/vOh+LQRC1iIsW3v+L830hTZ+XzWvYN0CVRVB0by89lrU0PN
IgZVBkveJ7FGZ0GWD+P5IQu9mLep93tlkioUJRiMZLghZzK2GqgQ8GNy8GLQPsyB
95XHZGM4eEuXhRsOKxt3YG4Q+KCiSyYE/sdegZS7IAX8w7jcuaGsdqMefMMC0JII
//hHC6UXnVryr3wRxjf85KYw/yor3JAKTKAOrnPdGxOQd9wEbEwxa3EDwvmriQwv
F9Br5WpV8e4p7AWwvn5avwSQuSD6Gglqamwi6G1d1+Oa6VT6hLg2wyEWW8sIEVzW
iXF0siJF0oxwUu1jcBjReuqwTGJRSDAXZYJ+jIoymdal79qz/rabAi32Rf5pY/p7
pvs6tIPh17fWQsvqyw5jBoEBTQFcxIMPfM0X0/0L7yOShPpGWi8Kq+8A/SQ+pZKJ
IK9dRwOvHqVHCMzY+vBd0BWxdrnxEZCYUr49gZMOpVzqAMiZl0iYOhg+HPEz00CM
mmWOk+iBDVvFUJIBxdNdTWbmNwP1QlTdbxEI4H/O2g0QBT9YRUlg5cXX/0XG390j
WjcxuhIJlfybVQS+IQnGm+XffAgLC3WjuLUtbJFxN1T5BrPrjyiupzPuJoNdWJBD
k6QnIejlgp5zvYHJ67cw1ZJgOBGHaM4z6qK3jcp2YmCUsxJ01+gYH/rQYd+MtsK9
Qy04nSn/6X+UIsuTGt2jZpLqz9jLRYywmERTO1A24cyL7m6yf7BrIpMYjCe18+ZV
iemic0PRrMm3M0JyTa4fb8J6X6xBViEfVPWsghSAgzkSy6PB0gs5vtKfsFJ3uj+E
RtjfbauKvNoFNSJLEby+e82RkebcfvtxsRCYJxx4DdaD38sj/kcH+1KEAKXhWIjh
TEW2HHTplex/hvEUiievWUm9ELP9L5eprukWvDLa1Xrb3nxmV6+sM2pMSXQxRADQ
JiQuVsXs0q9/H8/iktWOqrjw/Ui0CN4qw9NoqmLNMlvopCQoFgegCtR9NwEPbalI
s21Jzi/iQjLJhrDM3XAuBHgurZhr14O55ED9GbeYn1rFRyzEsqjAmAOp4cxrhdxt
lzcLlUcGpkDH/H78/oAYcUGg5u0g2tdg7jx5t7w9xkXyje2sJBLedL+689ihrmSt
nCRdT7q1mVGhDPAh/sd3Wf7IZohT+86IzTjgcs9lBhduBcRZIJ0qxtbAaMNXdJzb
ZtzUY7VueheT5wkiUVb9INAiX32qoO6+u0XetxwRlcr51aBKQCJh/ePOFBKccGcB
07sNPDFXoI2hp63TA2CjqQsfBkrtl6H5UAz6pAZCaOFQjPi/rctn9hdCCQU2Fevs
NnzTpvZAbMKMQyhv8d1uBwo52X8Vheda/prHHNh0IT7GCOd0jgfoYwHlzlXAEhyz
34nsNlR/NMl56DwQLcx+uP7Ih3hhAxrBd3XuJCa22Fc0OFnxt7NcGvRfvGAS/RU2
BP/fIOVl+YsQmOvh8HPKn+Lo8twnv9gnOQpPCCYMf0MA/RvJ0j7pT+jJKs6kEytl
pg6zh6cT2bt0sqBJaA7ztA+8eYxxfPdse/pfuUsAU7hC9vsBf7isRCiw6jqQEAcE
gXeuuua8a+j3BD+5j7OG5+Fn9BcBOipdqr94rgf6hGzuYaluvHhvV3caZP0Nkc+f
Yjdrgra9JdJQk/M1jDTqTWz8n0FDeCkdglKMdUVSA3tv1oiG15w7SZ4Ewz05S+iD
vdRHdVacrQzp9diVRaM7ukf/m3EO1h4pbrDbYto00fSOvRsy2omSmWXH/oKt3hyv
6tzQv4fuE+iMihMY3N3DDKBwrZS8Bm43cZdsz2dcTdF7TMQy1Sxtjm1XVJA+0sHL
FP8TyCNirLOUHXw343gbDDAhrO+ICbXq89l7qWP0J4F/q56er0lTHvYdzb1pp/lN
yWgGrv7nK4L4jzGMjy3BS6eP8CwGkP+9gEIFlvS/Cm5bujEqGKjVvEo8jfWWVS2/
f08ZZ+/GV8G2nkqPnimTrI18PQfbpqOE4X5awqcbiNvtzYIc1v1kGC0LyS+QU21L
dpkOXZLgmiz8wvmn4NM9FCc6JL2O1s7WPvtORcgh8C9tgqwAHzn/JPVH8UgbuFh3
OWsf+/KRMJ+5ovHncgyyM75oEbPk80dtamMwop+0ohRh9fDXdRTTU3tj0w5XFqGo
sDrQnbHZbh8xjVSjX8j9F3gL3Pfz+v/bGU6TCEMfbi9rnNxypIV5NCjdRIngg7Gm
/PyvtfS0bcLycwDjGWeRrbPbaXGP9B96I1Ren7t6314C5Zj7eZ3D0ZvNeFiH3+LW
cCR1kfbGwGdIPO0hd9xqNjDH8vRMq2hdfmZBF71h6UrImT/01uJPh0PNULWVRA3Q
xRflHX3GM36W1mQcYNambwhWJEtAScWLcdFeY/5Z5xYZh0IdbLrFVn2yZvnuhiB1
9kH0qlkY8P7vJgkNTV8Ov5K2VxlX9s3xSLRln7Q/cCW0jfuhnmUzKOw55SN0yLzG
xRzk1Vmnj+G6lIgROuneXGusPaJ49rzsxoCy/FkfLwTPdXk2j84CTr8/YnKKUals
oGqY/QVceefD2aHbWxTIXvpOQxq2w+kfjkbGdiFaweKPg0hbokLt0S8XWq8zqIoL
oCFj/FFTlJffAajTs1We02khHis8JJQpCx2ZlH1I1Sd7p817Jn+hBwaHY4TcqU6o
EQgZ3FNKiNLGgy80LbVO14lz05Ie5RuldqotCxvQSEpOQNP7BtgtMXemJR4KCSCr
9LYsxd92b+DmaAWNIEzEueZwHOctgC5LyOhm53/LkEtPBXzxYA2mdNEuB1zVPr1q
x50tVbGf17GXuYtV+RvguQnBbGODMoJCJ/a3fqQuRy7Q+9c7QSG9EiDhS4r1OQ8S
hrXk/rQDWEjmvaYNrTIfFtxfeUJUGNP73LDFBlBzEQ3GWAKmuiz57V7IpHp/pb7/
FEEXzy5pvIvDMyy4HCkas1zsHkeqtRVjhEH7+HSPjz9/JPSPt3Uu0pCru4+NG4QA
dYnRubYZcJ/Ns5n5dE6wv2nC3fn3EEOSr1R7iIxJvDPWwFu0ePdxtSQiWtqwVj+t
bbZsQfsTg+OZM7YRjSASlvgk08WbX96adG15U6J4DASFOfHtu1ZxkkOUUovXvWuX
FuB0xR/zvEF1vH8G1/ypuLBqIdhLXGmstHPCiv7bIcYdUjzPHy5udgfeN5jkjccy
wWSMAhoKnrCb293GofYXbI9q6TW8Xym1zmeC7RnU5aUC6e738f2wy2F2Rh06wi0E
v6IUd2MQ36LywfrCdPqsyebXW+CYl+hkwVXzvqkPGx+ZoMyxcwg3i6Tq2mlpLlYy
I9SIh+mjspGOkTzfsw6CGq5OBawW73n5z/kSRc1tPVZhPgE7TKC3z3wlQTD5PYzm
4QGF9atxZlG2vLYrWrWclFcoFvEn/aGb56aAJur9jOH8LQjEAECypp5tJm4ssWz/
gR6p4qowZkFo8M4QZ0iith/PgMJGn6jtHLUAoKta/1w8m5ZBb2pU7vFjF9JxUAeX
/N8wTAeR/UIaegGhgJ0oN8GlY+LZ1aFkkU/SVXBbZOu2q6Pc8IUyEAktSMwGqU8S
7ROGWMIzJ0YIkL+QUrySC5TMrFkBITXV/UOb6Ic1wZ1vUFf5T+qUkMz2K160sIM9
4/dk9AutU/JnZYruHSyBKudmFtNV1pTf3t0IgKe0VM2IwUPoCwVMKcRnCrbznf3x
PP0l2Ym5XZaSWwEwNm16+5nWnZ3b0nOik/4nFn+46zE8OQSF3Vt3ZWv4wxuyhwdr
JL0QBLmTs4JeZ0t7RdbCkutSvtuuAx+k2z7Mtp9CeNccRP6tfCvmwzMHOM/QVBpO
RhkgjvPrUJiT0hglV+XrbpCBJpEjJgG3oEfTgA+zXWpUn+ZA04JUakcMxnDUCLKl
qUB9Hq749YxU/c4Wgj7ojTOpyU5bYO0/LrUeNwc4OogiJmEPT60tmlQA/dFygbJF
QfCAiC8C4yVhX4kCOtKNtzd+C+wWbi3UQJO/RGCi+wcM++aVtS29wo/TMmXLBWVI
vCU2vm6zaH/vAcS7X5M5E8KhE20LWCjxa+jtBi8dvL3c05K8V2YwrMKcURmnNYCd
KuFzFc58S4EwGl56zA3DpblNPsiZuuInkd3DFxL9gkVec2YaXCD8jgEoFyt+h9kJ
dEH54CaiwkseAe/tSzO/rwBwCC4hSnRodlSkuH9o9AxoXD1Hv67AJWOakwineu7N
biBVrAmV0Qe+GhsJHLc/8xvF5NDNfrH93LSE/9DS4tdh70sHAcQOaA057F7HHBKZ
XrnyNw9fbRf9EWbGEgWjOKFyfvf9A2PsX5XEnh30xPF0a8gDipt0KkL0jdqU5FnD
zmoWphU4smPSFFb6fKcUQJedI0UB8L2BoW7ZvfQsFB4Wafr/cOP1pq942mLx41Z7
QLV9jvrPa7SAaXWYMGZnccaSPOM6mTB2alTtNZ3tFTmNRXpo8vYFQG1CI3J6vJyc
my0dXaDzGPjxt/EEB5S6i63lzP8iNqT1fOlqarF3xlwZBxJPB4XM1RGd97rE8ttn
uk3qLgfUWKYPrYkJcFcqEuMMLmugyu8xJiHPeluehFLTTuGFSMUgWPIAfWP18eNp
7WLqsQSwdkJTtF0QaAJ4EbGT3jL4PR/nV5/+LVDc6L8yMjueGcQYs1RP54Ri89/3
bW2b1EIe/OXEUwnovtw5TsGuaPk5Pb48mZJwpkqKDaUvKipcSTOjKANYFAy2mpbe
sDCZVL4upGRK2WlRxTh3vQ1DvDyQ2wvMzgZ/Ujfcoypd6dpaoJDhW2WZf6+iZWhc
XEdXbqChRU70lBVKHcxjgCOiy9VM3k+fgD9YbfJQZ3rx0I0j501wFdK8wah3fSDv
RAkP2LesWMS4EjHJCQAYNCvZm1sD0Jyu1CLJsVotqAALszGp6lP4U/BN5gSMl4Q0
RWWF/HrW0egoXmtaNqbYgW2qiBef/9r+qt1o12uX1XcM/sqAdGQxX0BJ3iiEFtCS
TBPX+rKzfd3nXm7rpon4lGXAqCHHIZgYZY7depYdCG4l9tR6P9bKTmSVVjMAQfKw
cnGZYFAiL58F3+oYwe/Xcnv5UEvYvx6KLPhNvqhALzYx9WLTb+kIrOoCR8xqGjl2
C6POzzxf40UelmZr2eXJ9YnWhmEhKQOiWhOFhRU5zPw+NfPMSwQ/7zzoXxaXReI3
pW2pXG25J1MAhwWU6YloSj517DBgFSrCeaUrcOrqsguEN0QXWCAMmfd66uaKbfVv
8sEJP4ShzYMcAjJEA6FnXj9utQXc5elPLjf2OZMZu9Bqx7GVeEkmSt+zXIa+lrhw
zrxWw0aFh2uLJUSUWeMx3Dwd/y2A50gFGM2ji89PpQn0EYEXXvaF/0yA9Mezir/r
G3PpRb/W+w019SB1TfEwXXQJD1wChvgavzn9SvAGmR0IT9pQHI2vUKWfG/D6Zt9n
iT1725mezqDF/vTHXr9lQWzwIogDUADYc/ISjhDXD1TeljXCZF6wHKfmAY8yCyGD
3l7UI001KMGtQpH2cL0eW6oEpt/V3UJapntBz9eMwuhE296BMsFd4zRGT74WxbHK
gKHE/95jxkN51wG7iPq5hnREejZk0dNbyvzvwkIdpjgozrUo17G4n4DEZPCgSTLb
9A0tTRjy3ZkhdyZPswzTiYoHJrk+7guJIa7oCaUJFvHGcknPO0HFS28ZKF7ZXibr
t//Pvfeo3eiHKqWY3ZF5IvxdBwL4xP0tGd2Myj+KcWdBQEAEOh9IEFMNzsBRrcF8
gyZf6pFl35m7TLatazhhG42V5BtvlsOI1cR/L9fT6TZk32DlMj07wAwQHqpplCjb
pzG3kepu/RJpOu75M+odcB26inh22CsfYTFwI6WIMd4p20Y8HhqnY1mJ0sm6KV2o
+SB+NwfyPofaSTKd4lAbTJ8GB1e6nst/Wr2sp16vfxAHAuMguuRVEGQb8GVMnlNh
`pragma protect end_protected

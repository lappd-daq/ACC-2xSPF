// Copyright (C) 2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std
// ALTERA_TIMESTAMP:Thu Sep 13 06:32:37 PDT 2018
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
AtOYYDbegVosI7bYK9YzpX9N9fQ5ZbiGHnXbtiQI9EI4Z+msFN1u+kxXDNbI0zwP
GOGFT0MNnkv6GhB5XYlDnqJlxnulm+7XtnjjVC59VJxy4G4wPk22fpdvluKN88g5
X7iZqlFI829iEf89PO7graPC3LhvbzxaHCVmeCgALJQ=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 12432)
qFVn2ZP6QCL0uRsmkP7EKWJHT1BeS/3g7HXQfMGkYyn/xKvIsolzUV8/dQOtbXrv
JOcu588Dq0GSqpwC77BlfJ9sAlJgdCM/fqif+GnCObKV0qQKnoPHfjuI+UM2uukH
7dAGvaJg6KVe2Ad8fk/Qx0196uDjTg6wrNZuPLCPCIFEQlHeaPziu7lHJBI7dWTr
2vpx4dtKmTwWxDse7anqu4STt/+Vf81vdagzzFNTMqbOb5umbjnc2K7JimOA0zOl
NpsQ42sSvL3aBBRkHPzImYR1AoEV2wjk4rvT5cOnN0HwjC+fBSSSfb0L6CwU8qGd
BsPXDYj/61bvv4yc1eOuy+pjbvB3CT2pdKBs6hiH25nHAgpwOFmCcl0CrLwjbztC
huVh2Q9gZ0Zc12VE1kPdKlGN8gYTGhjaIi79NAHj11+l3Y81AwZ47cjkFcku+iZf
u5nvw3eIC4nyOdIfdlpfBpVTC9/jmqYwjcmfI0vgcD++nX/vKaj2K7EixfJ0udK7
xeHfNWEGqYOgtymlJYaFbCaIIO3Fbm7qhbRQDZcY6AaPeC09pFOfHudgxYgIxnwZ
3uM6tK0Znbu0WddZkreRwSdA6KQ1ZOPwToQn/OQAYW+SBegfCu/1N0s3zZ9Wrfjw
UHzfe53qEqfV8EcPrg9EflGQhbRfb9uYjVK5i9PrdQ1sb2HnaYxCdo4ml3P78xi5
6EppWMJaHANjYpiw/lAUc4SCBRzfwjrrWnqF8/WaIBd5eJcl6n+0O7p66AHPxJp9
1xIiAxYnIE33vlRuoQ8XcOMjk1YD7ac8OxFlBD7SQf/4bbK6pUaoqXrGy9HaYjLr
SdDgHy9kQaNX/3tdthIwTDdHNwxg7+lq/A/+59qaLuffhSxbPYKmloIHRR4uIBmY
JqbGTAsZIBYC9knkK3G2bosQWRHWR1tWBmW1mi6hGMKx4zLXA5Y7ZxFDAbVLe1ep
1JtqaUHPrBXZ7b+0PD40xy/FyQHGWR0K66ZEADUJWmEeQeXItTC52Zt6hkCahjXv
N+XqrHyVWkryM0/A4Q4rT1pRYmav1lrhuk3l3vIbUmNo9fzfUC9HiXNSB3rJAP5t
SvNyVdaih5NkfYnYwbVK+Mjm2pKS/nos8VwnjKi3InOyKQmqCSp1k+SXX/441iEe
fmB3BI92EomKZ8CH7vQFjD0aygyoxUWGVrcKd/iwgMCH40YTkWHFP5+zwLjTzFiy
hk7TJ9/nufOBBVpL2e/TlZ8Z1Kl441cweAVpjQMimU4gLRJNuKo0qpxr5A6VjTmn
Gpt9YDP5GuVEUDCJY0IfCFZhQo3GN8q/f99NLrkyYsFdkIyxjqLplTrvFNdN3OeV
hB1WAeZ63ZcxXAk2qgfpzi7Mq9ZFM+y+KZwGI/jc8ORqRnOCbjzHwQR6SHJlRJJ0
b9/hG3b/KO7Yi7IHyvmLamIm+5WHVL+wQuONKOsqIjeHi1bxZtKGoqPQTDPr0948
pMK4mpmCapYCc1cpJT9Pywhjk+vE0QQbBGS6s57vrw8kijhu8AXDQvhUrQTasgY2
RWRrS7MHYS1iCTky2Z/CgZ0IxLN/K74u2e4e78OTVhyE06zekNcUaIJylQgcy398
juf50lVLjyaLrucWu3w/ERYWR8DzXUfd1zwoN5mzeY/ibKjLlWkfQ7/OHjgNMM2D
kDQ4pTyzOIYr5Vn2BqEjMfC0/1tOnMl9fJ7xNWuL1MQtj0a1y+TJH8b3R4rROdag
lE3FPkEpBJsPYKSd4yVTWDMwgwUdPnivKF/PpjdFOPaUp4eoYU85/CpZOC+6JyNu
f40cslA263jEe48ZST5fNUGVi3glyeNk6fkMp8pGOVgeCEvaVLQ73f+lenyz2AjH
bIk5+LsDYCPYLga8eJEkQtdGcz/rgR6abPzsryYFK64En6MuHDY0Qbhuk5SCT2CK
b9uUtT1m/+zWhSIZipJ+o21ITWvwYOK1FM5MrNelIN17Uunoj3dJmmI5rQrB8vpX
DzulW3FBUvpGht359J2Ku1StZ5h/tAa75URgwSv+UHD+fdQ9McXMYYTOW9vHbivw
jAVK//D9CrDyvjFiL2M0tpxopZKCaO7acjDcKsiOGPGmpOCh/kaHAR4SYcqtj91g
4hmm4zGqgcwjQH7DGQgIMxmMtRLw+bVR28wgIFQBomG2udqlOOLBpREMzJ+awyS7
QSa+Echel3lBjOkk6roKj4dZhxrJe5yFic7zQ2uRHMEyoU3KhJdleBKk8aPwt8Vm
WcXqZ0LdcojiFzkubZ4dNcdm+Qiv7LYJ7o7ZXWPf6cgWTQfg/uoEocl3AbVLsY+p
CWK6DtjXd5okjkwqEykNQZ6+OAuZPgjqHrrtFytD/tSJO6ro5d9xZmf/QF1AQ2eZ
jFC6Op9nIzfgrtcSz/oKZAjILM02htvMAx2EqJoZogXci1VJASeIDW6CeRr9pKrn
uwz23s4eFDrd3or7/bSoqiLV8WsSGcLx1WhrtGNFL0GjotErAE8DuwhvPRY3qTRS
7f9vgGh39dvVNOcTRV+m0DiUc7rZqDspBGFkvd14Dp0Mu2adqkO42BOjW3cRBpzo
zmAOtN+eKuKZM8RFH6HQIqxM1NILu78hCrSpNj1XudirGnhekCh+eDXPeCYAdcWe
pBEMzprrWL5b6OXsKdEU56noj0MWbzDmmFuY7qiDyz3palBf/OQbCSaELzrRNiGj
tiC3kbAP6mz5fvu0/Gi0aeA3oLNzX/TgmkmEjy0Up/gFsq8XJJ16nMeEAxJs8VK1
RN46jRx2o0C/Ipl2LMUsvBSL/0fi01vDOXo7rPgc+klrlxFYhdgWE4AFgJoTHp6M
S+8ryUdD6Ry4c7AaEwV2UyWVUmGaNxhAsoOArwmf4/mKQj3i7k+YLYhnp6lJqPpZ
D+amhavCIcN7f2AbQVswsDImh3QkBO82VXBXjIdevCVH8IoVcsC02SG4bb8CS1SJ
AyPohs6Teqi08teg9FxBcwE+f1oxqVdVGLmJ/RpLsWDdZ2wP2fmq9Mfxz2Vb/3pi
3GQTI+KRwuh+XcsFAuqEoVfM4IR2zcq6N/y9Mol2m0I0oH19kTXt4MpV5vPvtAsU
sKL49QvLqLlwVgXiFcrodwmXHxW2BFq3yS4gWKXsyUs7rP7jxhc9g/MobwILCgRF
VFPVJo1iPLhvEuVwInSuaGbiBImYofALRUdy54BpP2/6KKkRKmWQKhlLLL3Cpk6L
mt9hC3ZTrfMqg+ovicQH1bliGqehhgD+GDYLwdYqNgsEaWV7noPBaQOrmpqIDAQj
AXN56FuR3cd7vXKJkKKH45xcEyQD+ii9KWRD0DWdlnL/kfEmlpw5UjpoND1Br2JR
i11B9FWjggXdg5OWpKxQ3QZ2AVLan/hc2Y4/i2/ELpV9mrgaA1i59k2WEXbnDJfb
0to2LAygLmVvokgFmeA3LL+zEsRnMsqDWl5McyzNLuFHtfLBMmtVnSNCKhDRRBnR
nYD6yxL+AHxhK6B25GvxKtsD0xixtqSUaKG3zr9nXWAAbyyyaNow9Iwp8qt7/Wbk
QrrAnSBziJ9uGFZp2/TQNxaFry7ZA3L30DWcEe99DsmGQUwH22U+2DOaUtDShec2
+DygRvjeNb68OOa9Mzhwc1ZdgH4DakU5DCN6ClSn3a+CObt6RrpAr/QlbzCUgTI9
IAUHSd4Y0d3jS9/MLOFui1vUKrOIBbHsCp5y6SL9OYCnDvyWfcWIdZThs9ln+WuJ
J9x398/pWL/WgoAblZtN1m3SaxJ4J2c3FW7ZAAvUHYEr5SboQdVrpT++5jzppvYe
DvJLdb8/pk9dSpqN2WP61sZ2bQWj51mQZyZ9od4dgCksq0nnEqqjfg5EM3MOHLYu
SbeK3qR/aL10EZSLw+/3aUCuuPBjj6uhRSSXh3pQTeSwg6aayQU2V0Z3E5wAqIEm
s66KlXsQC4H+UTgiqvyYbD3yU3n4qbQtrVzehMM6Vk3QHCBelqTDTVqf2Xp+cp6/
F/Bt214BetDT+gTD3JYuEtG7L8KZvlRFH22bi0iSVtx214dy8fiJa9TMadUqaN6W
PWrvpFaVDigpZ4xpogR0HrmbEQF1MnjPDqHqkXfFixqHgQKbAJcx0uaJBm3BPMHx
oVTixQSaX3malmMUeLtcsns0iHrTbFxQ6tShsFqxxTY71WlP/g33AGaCX6dir+WQ
sXkGkWQY7uBTHGdQ8jOVkndfy7qP/UobQJIto3icKe1No0dHCTlUXFHH5QDG0dlS
T1HeKm9pDxceSaf03kgUJzNIAtJhL5TAYlX2sFXbuGDC+o2GWNLTh5LHRDo8Verh
+JCew9eMyrqDqbssnjyr/A0rg4400epSYqIgfWvvli1BXrT+kXcjS1FWmY7wmgw3
iEPSgSU2xE6oNFGAJcddqlhbpO5/IIgeRB8aI188m8Hk8aGlkghQrL2K5UMERcGm
kcY4OumcIDFWDTpbOthmFSp2AytcRg0EtOHPKCgiaeqkVUsjF+YI/3iLcXBQj1uF
kiZgHReXxp+1Jz/tADjtXMLtOC/FsHDPCIEX7UHRNUa7IAkElQ65dELeTJEohnb5
STs9v8cgdAB1D7kws1m8QTWtHOgxmY2pyHj30raUTX8Nfl7uGCf4RyHX3JXlE0wx
SHB63jr/o7YJUstMN7EThMO9dZIg8eo+ZsNU3t+yOk0NWy6ApIDzDnBguYHZLN8j
eqsGNXLwMgH99rbEchsfUmxTpfWQq91UIJfe/D/CfuIU12Fg+DfRHv7trF394y0p
86rzFYpEVKTe+Eov9QvGxbJZFNMW/eO54UR9cwskUTgDl4iFQdCFt+M6Sk3ERXXf
ilHvUXG/bZlQCPzjPJF7YgF/64FCpp3TFJ0oeVdxhlq4huYCFZaUvHCfMN2/yo2n
X3FNqJ8g/OpKyh2ZtrLZoRZ/yPpXL84H0SCrTAcsUbTOFrXwzNy6j00Fgh3qt+6F
1WkAJsMMQAdRNRDjkqRpJXO+vLb3aO2COlqu8swYda6+mHO+MdZUw1GBDrX1EZH9
Fe3H24DKS81JvuT9YLta/C23t7yGevKLXln7ZnkB3QGvE7SUJJVeC4IhKGvUgYQj
YqtVgsJY8g8UkJh8+Oo1smWYC8ICnD8YJS2j+NRSw5E7jf/1GSZraxTMHLWA0exV
erj2fCmPHCehJOMZb6Ut3Ya4fVYguvaYD/qCkDfwMYQihslk1Y5piCxcytjLHE1C
Fo95oTka2wzCwqyAVxw7paWCO2Ny6L27PLiAWY1ZHdUI/e/CcLpC5YfFZcxGFTmD
3Ks8oiJpsaFxEhgQY+ycQG96HJpEP18XnyqtV4sjWm+N6PmBQYcdgqY5mDKOOCTj
jwFowLr0JWl+i2ue/OjX6PqRm/18jPgRXD22o+CjEgCg2VqCygSrZncwiorZ/Q3G
2u2dfytpaDj6rpsApIW74mrBqynnqh8BvKUaXu/jTk8A1KmWw439efA6YykApdbh
zRXpLKoqOYR6U4UnTzTsH+wjrKwyZjGHmwi1H4kAWXrdk0X/6irZPmFe6xq4GMAA
aUWe5SsqXt1bOCZQdrxyWjJeEHU/CmKmgpWvlSs0DXjeAP9AQ1bhbcx6yB4xMnoW
f3T9w7+MDJeqQNOLfW840OqFJuGyHVvpTmRfV7UWTvNYwlss1moHOflgJ2mqHlAg
DwzRpvGHD10rtQRW4V4ZuG4f/njXe1jDEBRouhPw05FHTy9HFnW9FRJBCmKlf8wQ
vlm9026jzVCg/9NHjbi9EmsxreRCkdpjmnpn+z0Bculhbg4UDc4uyH+6o17vLEPK
ShaMZpLrCJMA6veqJTWcNgVpMPE/3k4HEmkYRhyN6RGsY6OR9WAp66klQa8/wdPP
opcgw1Nm8LsG0wQBy4iacTy0VDB7P6bHqvtlLCrxf1rZibHDYl2hv5L4szxrwsaA
NpIQswqW+mjqx1JWYBH0CW0In4LhdFJA0j72YLmWK0E/KJLVvZ5Pvb/kQVin4/gp
qwe1h5gXZL+ReCKtpP7L7R5pAWQGMUxYaPqwsGXin0R52wbnjOHwGLQ3SB/9jqs1
4NwKUXD2QEO+ybwiZm04SySvoRgLAhHrLpPZbaFimWPnQtFRyrIaYMbgp8UAcdEz
/wqe3egfoYtJ7MLi+tWysK/JgqlHzlbV9Rt4RTcLjTHqVy/hGeVEwTXntRyBAJv4
YBTra9tVn6vtXQ0LHPHhUihcmd3IeHYhjrm4i20sC83ZUcGNogti8BEAGPk9f3zo
knFYVqGFwj6HxvebozXlLzQP3fsFQAxEo6T/X0uyhtTm4GKra+PVRTaQdtdQz+Pb
AlD0zBIEP39rfzfIk1QGwZ5oKmFRqVY/PJygRUUv6TxDvS526Tmt+cZqi/Iqb0fT
cUKihFxjqngGqg5iwSfjTQJS56M/uEW0aELO5boTwIl0RiC/xeyWXWho71c72YSu
6jWqD1Q6Nd10IUzh/xZEcF1poM+DznftdiRd+Q3VePTMH80nx0cjyQCoq/PrABH9
WMvxKbqUwWaVsF/hXift7Scqkt6+eaGHlSE/T4PUxh/015iSVnDfk4yo0yLQ7O5N
xSY5+M4PS+KHVwyGcvSAymhHyhUlzdFrZf7XUxbab7dWc/V/mV+cyjDLczm4QEtC
LiJHJ4oRF252OyCSEQVCYNQqUkjkkdqkmpzXaRXYXmr93dScJdSupK4/9JKYjB2o
H5zgL31m+SOEtE4RYGUUS/rgbLeZXxlodWfpOpnMmoRQjmpdj3Q4klV3OeFG8f9o
mEDUYZJeuPQwlwWRn8KHiF6rjVIpFdZuzaGgggeEZqx6PiVPcJyzEs3+x3sQUIIS
quv9MfoL3Jh9SK1IeW7tb8ZSGdPoOBtPWDP5E+HKl2emUCDhXDVsPikqxEEF+Fe2
k7SiLWV40O1dteEUzjIO/vjH4+eqQQNSTp/WZwOZM4hNq75gyuDfEzW7WkjuSSXO
e+jCej4ukPbZ2iydaKbhYnHXHf3pQSkU9o4C20hvJdfVy7WmLjK9FQSNEWpRMkMn
AJW/dZ+psWaNv9rWVJDAfD1JV9e27sRNE45bNFCOgr6MnaYVFhsuFR9wdomA34GM
ow9QOAMxhDAS//CKltBFXBC8OB2/fTIFjMNo8+J+7shcS5wiBT0/c8ndMYBPyJ0P
I9JGyHHCSIk1Wk0EdcsduLWD2cV04Nw0XOLyNCTXSjohF59oQIEZI02JWomNggRU
UsfYrfUbZUdrdTb76SXCMPkrhohJR9hJk8HdPqxnkU99OB/H62e3bvydkIzcJmGG
UdB/u7TXpq6qu8E3DM753uRJmIKkRJp01aAN2wvJku8GbtFCulDtHJGSO66BxN/1
aIIbo8RrWJOcwtmc8iaXLoeNnA2QKsh1ifEEb5LHUfcZaEgWq6cRPm1fyFfaPUqt
vmqUyTH0ANHJHnQ5YO4CTRxBQG/X3cqgdccgCSw8y2+xvjmaXrMB1N6xdUQsbBc8
+B++BgYlGNZZt2npZ1rQfn7orMFbeRg1Ccjh/j9SX0uHWsTHcpN979G77r3hDj8U
UmJhNZ9+bVwmNv2kHLwAUmAXdOHUmCxpOTOmUiRdtbTq704I8AqNq2ke+gskVMxA
Avhy0fCNdFkxEOf7yvWxx7XcTAQzGDJ/5kVu47QShbK8pOse7UJiSmCjD/5mbhir
XjWZxPaRUhT+PrLI73G6pC327wKLUpDVBxdWoOCHyv2U555AgoyNZ6SJ3LtBADZS
u0y0NCytbzsQw0BrRFmNTwCRJ4A85dYKZrFn9TkniKGLryobudRTbh9ZuVZNRMwl
Bf7Szrs3C67ArO9fiWUpCQgyxj9kTOveTuWF4l1yhx7ZLaY7Wje/Ysa9DHrVOL7e
Db6kf5ialjGZUWYkxM+PQdWiXmujMoENYorXD2lB76rrF9cMr6GyWvxU2gXZnDZu
VjW8Y4kBiBPH3beoD2BXce9TJiqmhIGXOq03gUP1Rj1kNv0y6PI9tnrsHzbigqKw
i/Ek2ujxjWfI45+JqT12c3s2y3SsQY3Q/0TUPq8eqfM8pXOOKXEnOgGNEKpGDqt5
iVuqrnW6wW5WNXzANQTzy+AIFacjB7C6qN0swWOrFzQ1WpkTi48pO7mk0djqrsWU
Jo0dAzj3IiQXsj3QEq0PNmiC3aRi9T38EOa1HSp++88UdMYFJ4sQX55J1l4wxWw6
KTkmANqIreEDOghInEYoPb966T7uiZHuFHePrDvHu06NcF8wYy0ObLUO8HMondop
nzLYd4Q4rFzyMUnc4MwVCASbziAG+2W7Ss40GTuQXpOQUptt1wlhkmugTMxr2gAq
TyD2F0S/NR/e6UvRGY3kqZrzwE5UDB33qoRWoOp0WLnpm7TjpJ0na6MTdzhQDBuI
VMP2gT3WuO+ELnafsyloMB8ognwOntjk/0TNBwtq95Pv2IpZxW+vCv5+LxzVFd9g
3RG4EAHPPio+GQH+1062i4y/n8+tW62bxk6yQrYpey0Rkx4KkTODdSRK0pfenObL
Pm7UEOmf6fzx339JeAPm5yeDj1WvumP/cCMoRNt5MbZJjwiqNT5QJjNDSuEGP4PD
B0Qx48VtGkMfk38pWCxD6swTdpvyusRHAd8gKw0YvGSK01/7aI61Kdm/7oWXYkfM
ly0p6T2d07laTtijk+fqkUizd/tsGtKgLpVTM8RhrMpw0Qs4gUiEvN9ZP38Mbncy
YrTLcFGl0WRiASRh3kCJf3yqtsg+B36dw14LrIrXIlvkCxx9OQCQAcuovisjI6oJ
djGwgR4vk6zNK0wZvUvgLO//aWOWMIj/x4CHKel8Crkmx4VdOoap/KR9V9HEsZ72
kMwUcbS7iK+swwQq2STzeQ/I/DRKjqdQwrVHe9OU/U1r3YNCXoeC0WIncJASVfWZ
seG4lS9pzYHDvPfHuJAlazQJpKfG9TYTdduxGQOVg8HPRRVDv30mguZLZ26s7zDu
15k8NPJznE3/vAnLHVJyVxKKAnRyqI7uwVJc4uNwH9cPpyC37FNh2B2WMHMA0D0T
U7Zgydib6b+T0crBzZ9za+4JnpJqfT6MaABKQebYQrEERqv/gzFlQAAQFBIia7s9
FSMNeQjoAm1oTwyZ14MrO3D8EM90LYuKx7RzIeOKISY2GyBkFM2+Ns+7WSrfLHOa
DiJRnqPB3ED8L75jD/FMIRyI4tot57T0cQNkU3QWGXmN6scPekwIJss/6FIjHXKW
Ym3duRTThVgO73UwfFkO9CbYWLCZgl0h6iy8cfq1faY2nClbExK5/Gug1yfZLZQV
ElWJkzTe9gGsPvX1NoO7CtuFAn5TuXMDFPcTStsEpLgYC63VKX3F4wIzNvbg2FlT
vbBrzMbIGU6v5/CbLS0Cs0mYQuE06SG2tEr0Ggbiy8wsc5fOkQBa7CvWPk4XwU7V
YvuBQYSWWYt0VFXBgYYippx6IunoVBhLtKf7JUasS1iKSZzKAxm8f3jcWV3mhfbV
XiHnRr8jPG8j6YsarAzUt9A8YagTdV8MtZ6nIzeb2tmKeHKt+w0BlUKHwb1kcJDS
7fe3sKrhPQH0rCM/e6Y3PbmsYPl5+SD9jrjUKN0KKNyfk5GxX/Wa3GZWkbWakRlQ
Ayeh/Y4+cp3cKdNn1DEPJ9PFBsBqsK7UO94g7xl4b9YEi/kxoA5ecQqvjY6WEFF0
j/fus2EEPEY78loB204FbRLDnk84KnXvRihqED8ZoM9E2A8SpMgjt5OeFqaTESrZ
zodY9VzQ51I4/40GIbCvu7TWK1yCCM7RktwDzdukP75J2EDk8+az63w9kv5Fr4YU
I0QYan3P8im64gKTdGnMvsdrv9DE4D2O9lq4Gqq3Zr/03/8gnOMgiedEeLSORJ10
q8LQIZqAXUe7tYv4F33e0j6WOOJ0Kefjx+Jsb56c+G3fLHR1e15XyysGyANlB/vm
15Mmq3iqweeGbXnlixU+yqMJ5/leHFyS8+kI4xdDs0ExqJamzJsvTA8dQaFwvQBV
486nTPRTNctwrw97J4mRTyYAHgFXCXZbYmbGUggXwtXvc2ZbTvEy9vzDGjFs0URq
gV5raFWUq6A9niN0TnwIJ8uz6pLIryuSQKkv66P50rcNXnH4GRAoJbdcMEq9yB4d
sUaGf8N7G7aZ1R1N6vcqsQfmx1pmt1tL4u8ctslN060T45HFbnsyCt29Gx8/fS63
Qg4BXxcKOOxknhhYkGVl8YdtWhmhzfjIuqKn/bH/7Dxjce4hJ4M4WRRnhB1N2tpV
gWTOHfa045IiqFS0Qpw/ZJMH2d4TBaqgdEULb6SWz/3Vddi7AJ7dNoP/yxCU5ExG
fO2m9ndCfiC9fB7NIlzPWfRvVnwKxshBSyAvtXyMRMhAv8jftJaA8LVwRTyq7PUf
zxlH2ByKNkLoOy11BGds0oDasHD/nIvO7FBb7SUSkCcb3wIi5XjlSHDrs+yZjT+F
iwBmvycZDNPSdTrF7xFdvYsL6Xs79Jc7dUYXUe+M7p4UrmOAfqf9QoZKNIzoOd1J
1WkyHj59Ar2LjnTjkFrHfz0wC+3oVQB7EmCq/TYW23hUYm+K+jIr+gryf9jLcxfz
3s63B3BxuTUToPGnTC/waRxxlTFtPNP6MyTTdhYk61gFLDr4iWvHQHckyGvTHvMr
WoVq2wROIwMBsp/MDG6mU/rm2TfHT4gaexLwWKxyYgLIIyM5fsPXzOYlzrbgCbZ+
OvLUgZFQriA8E8oCvaNEVObN6SXB2JBellsktnZvK6MIykPfdB3I4NFsYET2rCsb
CND8W3/31/wzfOfQXZGvejf+ZLguNtujESFD4MDd6R+5uVj6KHXNI6VtUhLuKQBy
nh5H4LO+TYheOqprVmRsBjlRs6HSxpzlZQ3nzVBt5I0xVH3QuYpTpiWK1z4mG9Zb
KB6MTEfIYfPO1M5uR/JnoBYqSgRf/ht6M55or/Tv3waE9SB1Y22RM2dNHej5Ua57
xUfpWnL00pZTYpRHMuDWE4YiLHQ3Vu6kuQIGNzMA0B2vtLhCxHBDXrKsJtgya0eW
dvxT6Y1dKX4JvNFbTb9QHpvBEzXmIInWTJfU0mI/PPgehJWLIfwC/rs/8Q9kDpxV
QFFeB1fl51ZWd6HI/6xVIZEcbfOlClNrOlxLVdwfE8mnO3aBhg3J+IUY+Fxpkurg
tqLO6rBT790wUwgqEKev/uf0QTIGKRx/XNvD2eonCWAxiUtgkTpVSUO+QUscFwE/
XJkxAzFledeQwipenv9Zn+TfIoO/Vw13OmeDo47RiLz/e+tNKTEUIPye3JTXp/FY
H8xx7QX2WwxiWVYpnS0pTLKgt2IjNi9LjiDeWWkrdszjKMyBEgTgdKtD/a70WsX7
sRINiDuPDVxZuMp7WM9RRgDlSSa0/dGTWLMtR8h6UOYnCoQBQzkWMYeFhKCb766k
bXWccbBzdMPrdUJH/a5espvJgr/fvCs/8sdKZ5Mn9oGj/aqXvhBVBQ3SR3dRq1Eh
5JcB3iENtCrA6HcEyBHip0b/djAAuLNFyaZhaoYlGkwjg86sKGuk0ACn611KtuBi
QHN6O8GAICgHfTn+Cn/VTIE69SBYZyEj8TN5DKWM3yn8yaFtLis9SVLkbvmVWmxj
gdiltx0gGMA/Ae+KSb20NQNR8ApQTjMJF2PK7qoMDOaiwbS87vkUFlB3SxDFBND1
zf/Yf4NLKyUq13tHcU6Q5nmo/UXJNUFXZ2bH++ThbggynPD7w4KUXOj4/c/Xkngy
lS4bFVXuSW6AKuMYfRws6o6DalbnLQofzz7xBMaPcJl5rBQv0JJfRCLymfiCruMn
cYci86HLo0134PsXzHG/mQHtSrsSF0rheFatUUI6ooTtv6mZf8o6QDShtupGUh6d
531qRCbxNq/n0+a/DmKpGAgesb34lxGpb/MYUFb4bZVnY4XPRTYsjXEAcnPnSFMX
cR3znXhVj+W/izsW1KL7jhVBa8SDbCZt8IdktSYTFRmaX3uR5/bZpvWWE1Zvs8UB
QQrezloqb2I4SWiBUlOre2LHYoUXzaE3pj2jPj3yjQ3WYm+ZuPwNJ0hNNC26tWZa
LlGRoHHUN9BI0Is1XlVOxaz68VVki9Ilu4/50kObVd9y99VwWiuSUhoSN4pQnqZu
c/6137ZiO8sHw8o9A0eIUgvI8lLsJrClHTrAFEFZa7D9uIQ2D6cMffCSPpwMzMPm
ADyexBDOVyWC3ga1H6UTloWCzEmUQW1QhsoJMLy014BpZy6acpf+oIemUcD8URjU
9KaBYw5ForaG0RHFH6VdTYzo8o+Diy511vWm/R+hmqXqMvz8l1bE0XjmP/nNJc5U
oQD427oxWa60h1+e1bkhImvWGsUdBdz0UCTnJVz0HmOsze61JjS55tua6+m3bVOT
OvBl5CEk8209Q5KfiaiSIUcxb3+gbR/gPg/STmEE88rTK4i3T/85mFIWkCsc7SFV
VVLXzpVr7erM7l6flowUCOMAkPEvLBAH6ccA5CqRlIMzaKbyJe/vDe/TNZuh1RXP
/X5NVzYjIOaA2hMlA7lfWqpvHnCMatvca4470qh91CeNfCNI9MDi3AzRCAyxG8Dm
EAzGx8kbOZsT8th9JVejIjmN3gU6jBbHCYoUFYynzARa37XFiE7JsezY/QOl4eBI
iRwDECFMMwZMIwVZJgmebYRShtpu6Kj8IBO9eRIazHrpDnHoYCi+c1Ki3tSqO+qy
OD5mJkJ3c7hqB7UbrSwQnwp1rXj8dAamctnY07BAGUSTfas2zNFlrLvvuC159jAi
o2erQs8YSDED+Rx5gd0Y2DITRGqboqt9RgYLYREx5l8Ys4SNZq0MYP4lm+xzQr4J
50T9QxGNeoynWv1+Pl9w1pxSS7TgNp5ByGrVDJVCJxel/ZVa7s2laLv1DJQxfkkR
Tcbf7/UEjdMNPBPWUW6IH57IY+jrUh/1xxlYHYr41zok9uehRCOZ5m6n6N3yhpj+
u51NEMc+t0A5awr7aXSQvssV5Z2lTD+CO9cfDPA5HFL9HAY7drGLubOC7thR2zQD
LlKTWg/uMzEx3Sm9jqHjlGamUWkCU+pfoG1lbwlaq7iYnjMgbzm5JOzaQSMqveX0
wGHmuV1JQBHNNY9IjavKslW/zRhW+koWvO/ALWSxpWL9OqkYZzjiCPL5esDZOrT0
GULw0Mc9SmM0NTb8RnM9U0Y8wt0zpu9c2tF92r2M4luID3zDroX5TJyOvxZQmJgQ
4s3yosqDAXhtLqJZDUKbvY61B8JzPQqfK7sViAr2J9B67fzHEC+CLuEV5gtKq4By
WkiMdi2XCXnBgzTD/jCaCcTLkAOquqFga8RFQ23DI2B1OWYj4/Hm9w7gaZuhHIlP
2zz1T4gipwyrj+3tTRAc3chxP7jYvVoY+rexrNBuOlUm5WPZ9B2puFlNwqtDUf4Q
4Y9xRvY1HtluQECvDdvS2iIDpQBrNroJYX7ttc8gofHE6+Dvbmh4QVRo1q3IMmjY
B2pbsoSldCPdKP3HWMwZvb6BwtKvNQcyXdE2iZ5x3SygYxdimPxCnAS8UIMCNve3
OX3fK0Q4d6VkaW32ib6ryWQesBM7wBbYSMDvY+DeJ3iU0gk476JI1Rzc/guxPMxm
IT7ZMlbOjmvO+pO6MPrIIbfCL0tPfuJnkSoANJ9Y1jCmIcBnQTopxjaZnEnaO4Vp
dZrMknvO6CA6gPPgVaQTkYz8FQ6nLn4jzDo6PGW/q0vW3Wsg6CSKwYjTiekFmg2V
JY5UzPb66pnOjcwI4Ut/GoBPVRmrCdfk63AZEMTdHkBph+VGWBfZ8ej9pm+vLIof
iQCGowLzI4PnSO8+D06MaNyBGGmlBnMTMqPtTyYGWKPPmlY8leIV2YzRbL3V9fPs
I/F4WCAxszhgojk0Y0YNgMkiXvBSuNBPbdkk9NYJUuFpww2TyHy5lbZS8/QNyAgQ
qoXPGB/7GPkJOpXH4OH96Ipi/3lXAK9VCozB1pKcjo/rqRChuaaATbVBW6g3C6WT
NtCCxQwmo0CzlQF6ZEtGh6rSPsk1fFVM/+kzKnMcKQIrctLGdPYPKuKqlcZ7OgIF
CWrNogEUTkeDPrFFMsbU8Ce/c4v/GOW0DGHfyG17QvhYACFRdSo1GQPwJKoeMRGK
6OH9WahLECSzavySRiHRiGsZifugYsqArEOUNay6UYKJyYw+7LJeCo0+sDOvfBqZ
o+JDadMxgeSutpfKMrEORPy2aKcfc93MFSdToH8MzayeUZ0hyNwNJM1yndHFtYiL
UnrWcefA51FyySpnTOwuCpG5UC0h0N5PFhctdtDETdJ8kPRnxOHSAz8U1SZEJG+j
ZDipvaw4lqmpFXEtJJFYm/2NKpCdYPZAwPsqVITOdUjy7WtMDLdQvOxURmP5qwnq
ga8dIPwselxQ1PKKsgNzsofy3yHB4PpkNm7j0/Cl61f68+KEvC9vG2ievXyCEJtT
8H4F3LPEUhbNVtX1F8ORbFgvNRXj2bzGedhvwXaTb+IrRL1yrPz84V3dqFg5HhU7
sVBUOpTxwVV0bme0zbrlePkMjpbVa9qW0/vfZ7Pwa5fr32iaUdSbVzIDONPiiURE
Dqmu8wOowE6bImo6AQbo4LgeVQsBx4D1ieQL7hVuWZNkWlRUZoXsWC0U/TED0scl
fzhadQQ7e8pSgBthUdi5lrueqelMFhmavxHDKfDdXmoAmpuTe3a9OjojkTL1a0bv
OJDko7oJOkya1xmXJY13C75hHZVPfAqLw3k0QkQHhhh3baCYKaiL1PPxkAl1ab8o
LoDD+jS1SifZ7osAjZJUoOL1uB7+pD+R9e1dLD+ckqNXPNFOJ69XAZ4o+vuzwrhY
mz1bVarDYOhSwaDqq2250GAdunfHb7lP4jUZMuB6+XdNaSJAmG1trMTMZzOUKPko
Z2aq9StwXj9aq2ub9BarOcc3wAaJfG4B2T7ARIdE4AC/Pq740dtx/fO8tIHRFmNG
rIGGY8RSFxsczRKEQIGYl7XWIo+zjayyQnku760Fjzq6ZrwSiLO2DibhrEySFfaE
Nuj0xAYNooAksC33AsCPNiP+3tgxQUnTHM1aheYWhHutiRpSxRv9xwwdB18o5vxo
qbABgK/D15COwEmL0VHSERQO+5aBlzJaC04uwrZIpbqahwvwyXJ6bFz9BfwqCLIp
oDuFvuQ+c9736mtxdq79Fm1xsVMwY3r+yhKaYYE4Y/B2id90su+pKgq0gUiZpd5L
1yg4z9BjfVsRqsFip9KIhxP797KolzH3Ye85pmCQXIG915XE06aRRjWJY7GOcPwZ
Gk+cVQcVEoytPSp//iFlgXz56yIF8iJm3fEzKzE3NwTz98XYXhmYjuX24J8yzHeC
XqZm5PDp69uIRCCPJwtIypucPGn/L7HpUazQ7bmDgHVmO5C+dqTuKXjpoTzB8cHX
Gyet68LOCFQZ/R4MiB/26dS7ZYa2kZo8edMRTjKtFCgvO+g7cu8XDjYWxK+oDO+t
ALKrQKx1u2S8HZ69vYph/jIhnk0YYnObK1qrzMIMr84g+/4IHOJdBxIctYggYBTd
QcV3HfQrHuC9xx9czLVUf2HiblQZf+IAbmKRr0FiOK4VOtEab3hdov5iAGEU5WiG
N99gNp7i0DKF+YPXsrUaWG8oqelOxqUyfCS4JutwkqeajgtaIIhtbWH7Lt55hRhx
h9gHFZ35BCw7lpoYg1J69lAhRz/8CAORzIAoxAKXBeERSWLl7gC8rrlK4jdWwvxn
r4ZM+0paxG/T7Ybs5Ryk7ZeftAiK0y+9qxW2VlMGwQ0NGf+BxOGvF6Xs2FX+W33t
hQM0+nIeUZJFQ01oCtHDUh6Rlo9RrQPaVbvalkn0hvdLjZPKL+I3dDFI13usZ0yP
CAARIuwxhChWsJGtpzkdI4dXnPFlEm+4wJMhJzNFv06VPmTfwmQ/Lruy5mZkIQdx
zDYca0jvdoIWT1eooEoxYwjY2VIBYdmDZPn9f4C5CW++SayprpcHmtYi67IUt9ki
Q40feMlXRtFtqLj3VtFJMB7MIoE9TY2jp24S6Dv9CdaxBYcLS221KZmV87IWlNOS
8pckcnfezRM4uFmozKLoxs8fSWrlC/KMzvVZbFwGRzt3idlZ85K6JsshVf1S2pAm
1TAmjH0QDR9BZAwDleDUyl0h5ixJoLsREPOV+ibszDc1k4iTYRKD1qdSbTU6lyZb
jhkhXv0yCTsG53EN21Rkk/RtLKWSST2v/lvFGfaudDg0W84vdajVYPaOJvD9bFC4
DtOI2Ziu0LyOlayXiAqQuj72o2mkZ++yffGHgLeDcJo4WOTdG6TYwUUwTTW87sur
9zd1zq/3kO6we98YqrQyk0MTSlbpfnoYMJiZzvTlRP74+PHYJau5EYrlkIwGKgaB
GEZFLRhv5uoIsAuYAw6akv6Su9fcFOHL416zOCguvja+F5vxMj1VhumKCf3+g9uh
b7L7X05O3YeStkOEONNVUupqhUWn9dTHmk3Un+3EGUCYsEX29njG+6NsdkQuGXOK
VPhtCCvBNp5/iMtPOoK+6ib9s1+Of7i8XXfQoUK5mzCDJ+IJkXF0SE/zSftlJyHi
DSjON+XG2Wq7fAAROooCyT/OdsLj6qCF4pYOnxR0WYoNOmFOsHV0MWc/2k5L6HKh
ukk1evwsMQsWXDa4RsdubtnqshyD5W2hp/y6FoLUua0jDvVfSSXvt9y74y7mWI9r
`pragma protect end_protected

// Copyright (C) 2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std
// ALTERA_TIMESTAMP:Thu Sep 13 06:32:41 PDT 2018
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
QNRUSQK+qfBKSBKiof5Oe5BQQpJaAGLPEBPRiAiIoX15th83tXuItNYMgZ+i5Xmg
QRFD+JvU2Op9mSMppMzgpOWtAgzHhQLyZn9+skryfLOwuSwpp9co/u2NrTLoLv/+
thgaKERBPjQi3MO63+zOq6/huWrkS5UfdCKLdvlbRfk=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 3792)
//z3ScOIIQoWqpgwjrUZ2A1RnozPaKQLMcc5rc7RFIYoogd68/flE+cUE1BYaYVG
x/R6lJRzvbf47r+0+YyEfUfpohGfW0PnT5kEKdAQaZUYCOMiY4LTLfFDmWqgzjR1
PdcfSOUceBsF+Co9B865ZJZ6dNg/ExxaxtUz5V5zZgADoons8cy0/6IClazw2Auc
58nkr8DKNv4WWuBB0fFR0iz9WlDexkTPYhZzMeA3UaBvyfjUDk991rERAcG7gMJM
AV8VgWkmh3k+cRmhAU9i+OD52E3NIdhh/ZdQ+EMVyFw40L3cUANFG8F+f31+vo27
+xQ1gRqep/dB1XXr+kZZL2uNA+CBvzbHXnPIGO3hNLe5pBPDilC6OFwrW0lFpKM9
MYyiC+NaR6m4buJsjlIr2T+5XU+wB2KbHW/y0jyksRKEWQst+djnrbUeDpDpDjky
HY+anV5q2Qv2yf8d0E2b6oQfBTfv7kh/F9aBXzfcOrOQo+kyo2aYG6O4zPaN23k+
MNFneO/1dLN09wGY23dX4pPIhcp8lhDsGP4PuBlOl+R6JHwaEoMPGaridZxGj/tL
x0B8eVzL9ImqSJdqRksZKdQ0O3MduR+BRUtOsyrosjQAWqyUJirLkexN+pmUPist
6jUOplMxoYimsEP5fB/7MfTh4KjQmW17qMu1gcG33NwgKer/frD6H8kAGFisDE+G
mLc5wjoSLgpiegRDVQ4CaUyI8xEl/dE37RkWZqn5bh9Q3vTxe0MEaLtHDA961HfN
cBJJIFliVNLkUNMAHxhcJ6N3rmSVy23N2t/wrCXITqWeeQ5cICKz2mcr8czF+rpG
iDTUAwZVhMPwkUqorg1n4fodgQEzu94F5NQFnPsNenFFM7xPnUXMztkEhrNWgAQ7
zwF9e7aD8Ko9twL7PUVRvKiL/bcNhyEaxbnmlIbB4zMpEaHUM8a85O+deCuXj5r6
CarE0XVd9tqnDt1rBIR2ThMvmZjRzY4HuBw6gUuW0lFO0VEMA9OW2F6qS/6NuvSh
klW7JyAXvsNYysKFTESsDDlLVZcI0t6VlniC3xTGFwnsOmpxpSbEwErk08/Gq2Oh
aXLtpx3Z22glaEWO3EtXIBdoU+K8wmISvVuR1zSGlSnay/4bjNH96Qzn+Xy/tfZY
aO6rgyzvx0f7hB2os5ODdXnJ83w/Zn16YxPWJhqS8XeHJr6/GGr4rxpEZSGd3+4j
Bo9aRsHNME6ZFWFSNBKZa3S1wayv721ihB7oc6lTznv0vhhQXrh3BcFea/wDUWg/
gM00HD1UOIsctgSpbfcq+hJw926fx5UJapxN7+Zr0cTo0Yo409Y7Y0LN4wYJLNo2
wfNUnV4arlqjarL+ooP7eQ5+LoPjtaNfkV40xJK0IueoR/UOqchAuV3lI9EwQ0WZ
tlZWz72tIJ7C+HSzctadQASRgeggzXQwdEjJp6JqP3RzOpwJGg5JWZqrK3xZFHZR
OZGCr5Xwmo15INX0tFpIz7NUeI00Tw6lrzly4KdklK7AtKUboB3Zt8qPabdkxgoW
KASm+BGqYQlkUpyOH/FEOyyG39tdqO2uAiStbA/pNt0V91mEasr7B/ik7sfTltuv
i6DWUIMLgSRIPZWwG0DgYDgjxWFniNMhltVTVhFxwgw1LVnJGivOL4eWgMcQThvB
uTFl10OclCEtMm/TCpvGBlZVujTZyYvnURdJMs6z9xMt/Jhjpi2Zr9H04Y90Ig3n
KEWNg2wtSwEESlT7AJm5KdeBtm19o6KaWNcJDBa+7xFuLmw40267PN8sTQ7qJprr
Cr+R9f/saldxnPIFpZtEUSj7hEPRUJZqwicCsHhmRY+8/cl8IEQJGmLONHgSlZhK
veSlbAQHbCWtZo/+alMzHQZ/LzbY9KEx+ES1MV4JNKiWtSb83Uq3mYtIbFZPVCxl
mPWStJsOyKpH7MWlHlr4uvJACC9/iX7vQTohncO2COrtu/ndTP20QRPJ2+G0+pU4
yXLlMw8Aml26gbyka5GcZh99sUJWWOzytUh5eLthFeLJYltBLJLQDyddGuL5K6vf
LHnLjpsbsIBvWzQoSiJ+E5E2fSKkyF/4HQ9OGhZ45w93sY82ZiHHvEoe/tNQmDuQ
Z4ftEohECSMcxuRgJjwgyLpwtv+YnAdJLSYSLdB90VS3clXYuD8OKz/FcWH8tpLE
ub3aSLd5UZAp7u4zp+RsCua+VzHyyCQ89xShD7ZS24obwbm85kqb+Izvn30qG+9L
vXBzhxSGQ1Iktz652+zgRlp1tu2Y58+Zdpt9ZZZ4ht9T5WiqXlwg7xZ8sHrV4LED
ZLteW/UwmMPGoQiXGa/ioLKjCIZLynNy7jXhAov7bbxprR3pD/rtZM/vrZRFfOgI
pnBBim6VVP3/uQlEJn2zLejAbjhDtJETfxXcporU1AjAn1PrhFah7fEDRfjG+oIY
nPOx7CdIOB6p3F86FYuoX1LWiUMAyYsJnp3YqGR40pBldMfdwTv3AfB5FPQ9IlSU
Trr26d8pWyl6PbEwIzObAno5zZ1/b/YUOXfQ8wvDqlKwQzi4/vjgNuEBUpo82sIm
gjhJsNPFN0gzQlhCuTZJrGQz/2vT0kzbtuWd3XkdAVdWyVGJjjSnDp1QdaVVxVtr
f1o9DVMqZobKId7fBwbIvDZ1YWpvgBamXOWchaHcWfBIfkIjdyrQs9mdDRAl2rEP
ZPW7U3u9KlLeFcJFiTklgCfFGx1LGKJxOpvN8sKtqobJoOYIsO8dWoZ2d6dj4qe3
WamFZoMAI0GNFeNWl8Oc1mPnPt9xe4Ushs4mZ+WNPhCpOJcBbhVT2pGlwgZFQkqI
KoM9tWlUP5JdZEKfG67OQqDM/9TV1p8x2pIvsEGZmWzhV4MV1rgkvEl3AlF+/FYc
uyjPKmnKHKip7CqfcMAaUzu6CdU4IiW9CyBmXiF9cfuETyOJLHX94rueGh/GP6Yt
8M/Ogh3r3PehG+dg3iwgANIk7uH1cRRmZVNkV5uPgzZPP5mtCSbqsfXXw1Uar9Rv
IzuNtjE3MtKKTTQKIxZ2yidUgGOFabFCtfkBu0qRCuVLE6dR1S7oDeQFrmN6eL6D
RLabbRdZ/tcZud/t9gehwZVsCYBt81ujQDSJbVRiO72Ws7yZuaLcOhsQonVBi4Rp
lMnlnrYmopXr+hxHH6066dr6BI805iCPe2yhQY+5wlLHy5xSbINMutmjuKZr65Wa
1b3hdxK5zO7GjnpkKwz6gRlnmymBjYBy/CVw6HPkrm8EGDTSxlOIrLz8qhTjT4RS
sY5zGaRp1XC8/IU0nh0/IBNP69u0Gr2sJVqeZ0HqNfRS79+BRp/k9wXErp70CJWW
RRoAzMdYB55crCQq+ZI4CoHmkSR4CkPiO0NInVr4eVrryp8AehqsasXpOQBPox+u
RuJ9/mWd6e5wUuFOpFgLh5BE0HDqJfDBaQDo4Sd/eJ8caEwu8K78f4w6QFmypHYm
Tr2x4XvhVx/VDEUZAS0Mw1LYOQUM3RA7t3wRZP87wQGzXnvCLuDi61Esd06lbsaX
/YH5U8g7e3bFcdlnbaWAfWYLTccMUgXDrd0wWABr9uUYZ4tEyoBcHA2z7w66tRaC
yJSCo4HCyLWS3nEkjopLwwahiTDDyypaG1U3aCfUWQ+c8E2BUlaosukYnaivzcYN
9q6hL/K9ZFX6XYY9nJJocI9xShZ2a9ZMLbZfscJbkXVQR/RD5SF9+DSjBM5fG4oL
4eZNGomRuzMKuiTxrda2K1qcZXuTW4lS+6E81Re23VahTuZ63XKdqDENzWYcFj7v
7GqxWoHmnHUSUMZe/xx/hxLjU9m2lMGMbCVwzO556x09zZfDHkRgfmamBLWIISNy
Mmfs8qMPaeo7B7QEqlBgfDzT3N02sQ2119y7d5vyaFC2+93niZZqFAPnN7vgBz+I
qGZchf/gt+VFmgjB4BQ3PukQCSQp7h+AWwey84PFAoGGY7ETRxP5lza3nnhhplNv
Ci/qjajM7nXVYYUIEj4NYJcSzvW3ZfnjjiC30/OZQU7kSBBOfMdQgiZlISRoBLQ5
9bjrtt2zBBNn+Suu3ltBz64VJC4VV+S4dZoV0GTKO5pKJ+TmFd/kE8CVPBiLrCqS
elWCpNBcGmAi1R0fTDpkeXTLVS90bS2Li+xqhEgTfRUhGjMHUdz6Jdeo7PrNNFCG
5u91kfL8rAZYlHsHuGDVscK/zOXov/syWsdXWA1bHcG1m7+1wgfbieS3OG4ADp9/
NNdYdTNCjOAuKSbBZO94vMgVF8awpLsj6vyNuHWH+6ml8j5uurpjC17N50fw0kgF
3KkpwEn9zPTznZTYkTpC98lSo3a5PV7RjWIsF5s6jo1EoQoncapXeWYJIciHiVsV
T606BzPzWb7LSDq566hRhWkObrcXSRfvlhmIzmVUM+8Sk5hahFF4qr0DozmI3AZP
HgKUb86IXJPvHpQX9NFZifCNHjNj9SWmIQch9pwaHVbR9bTotLrUSPwkTaelV9tz
0xTLVGcnFE9RG1bIYc/0hb3SWzj55/jAg2Vzs09Z3C/VCbCv049N7qOZzgw22Vdd
teN7ZESOksVkR3M4kDBEipid5SgySDZw3EOBpCL+cDp8mtUbyNMNpaDTTjrTDvcG
YHJhZc6Tg4kLSrIgyejshuDZPk07mVOFEvga46NRMJCR/vKfZ4xkOmEYaml8ZY+l
+XzPpKGJK6kIZmsnjN8rsR/vI+hfEsJkWAF+cof7fW9/NfpopFPFHW01v4HaiWNA
afUdNbeUHJSAetDMDOb/yleOCBkZyDHjWNyQTdCwm+gxXTev/9Ue8T7AuNF1HNlR
XXrdWCyboL5ywEn1U9vyuK1mp32qAl2KoQDF7wnven7Sge3ib01JjyXye4Eya2ky
Z0v2/S/aLWVVd69cdpqvfvVgNIXkViztTfRONBVnMWvrLNiflMrmI8gSjzUPWsNp
KrtiZmBGB3KWcg/9RatTDt6OmkH/qCLiChKZHZ6BxG1AH9vnPRW8ao7e9s0CrhEk
pAW33c7rOQ8LILF7m7xhxmXUROQb73fw3tNaQEh6ri6loPMc9kozdhf8p2ZesWD4
`pragma protect end_protected

// Copyright (C) 2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std
// ALTERA_TIMESTAMP:Thu Sep 13 06:36:50 PDT 2018
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
l3AFY6nRpjPI1/S9c8G8RhQdkuvCwSxNXRjeAEkCWOMLE9UKHewMPX0xnb30eVvC
3SfK1EtojsIm0pNPNp9ayDSl3zsnPgm47Pn0/OThFtdKIN88WWwN2x4DtgcwEmsc
mhjhbUN0VaUrzoOKH53RaVCJZ2LqeD4qEE3xvBMZvfE=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 2224)
OsV5MN0pM3146U8TNcuxQf0yHNuf5YM6Pj6notFHiSnQfeWWqQOzgsXfO/nSAPgP
G/jPaMIMNrAn0BRAWquKeuAKXo8EslO3Q6aA5OktTJHfw0R7hDhNcjnUszZUsIT0
USOwllcBf04ws6XKuTQPlARHLm5EWr6glQU66VnYnyZKuO8FLVvjM1VekaQUYBiB
mHwW7Ybi2GZgRToR3qgnlb+yp5aXGlmq8838hsszmeWBE8u+XXbHVRLyS/jsWSl2
VRA1Spg9OLggeSWm32i1+UprOmzpbhdx8qtcCULLy+cNTgP6zYiL/3nO8N/NtjZe
RVXhgMpadF6KueQyB+Eo6YTqxp4rkVtz7c1pKf7rPHpqqm2zKxFBDkWXUmLy+js1
VKt0dKA/BrjyQ6creNqoef4Hxgyjr7du+MSEyPao04AOmDQ8PYr3XkYQXl0WkPw5
7587NZ/7hZbFQuvIngymQchrK5t1X5JR48U4M1bzhJIZNIezjUrUarPRlXXm1nKD
KoiCR+RjH5+YmCtIsy2DXf0guKI0jON/saT5g+xdMwwsA1z7pVrNheBhpvgn0WIS
A9ZL1dRGmUnOIk3RO/kzSyIhQMUSC+K/TijXQjF9tOfhIZaRPpcJzpvcAlk+bDvn
4AdaXcO3TsiaXFAOMG4e/188zhX4SANWPPzr845mVg6hIuBVoZAf02BAvVEATn3K
1GAOorsRt22cfcFxw3zzmhF8Cshl1sHt6xwFavZ09QVTtm2Pl9aOo/sAX+yKlnA1
dv7QCq+xFae+eVOdlicgDS6EimF3VMMtVFYu0fpoaUaW5oKRhlNROeb4DV71VrH2
lkR8BftlxzEypiHOvPEtW+veDG5qFVad3TYK1bq/dAFju8CD7Cs6pLnWKGQPwoTt
4IZk7mBP2tn2nTJbsNVfFo6ECOAVdRZ+eft+Dek3ZwE3LcHHHaLr8GQ1+ARjlaPZ
QxTC/WSQvHWyiNZW3edrI9Jv3wXNYL89Q3ioAUFKuursLPy58faRClwGuA9AEU+e
6veZY6YBYtzoIUwYj4p6sLjeinky4TpBXsalda73Qjf0neqi+Ix6+FHeSLkkN4nA
7a2nXrQUrdTVASUfGuZ1ayLq69vWHbchEB8UCR9Qhb9b5+ZTWpis+ndwd5i4o3w5
m0gS/JwDUGHiiSpeZ/q9BNILZBCVLiGHF8zHSNGC/E+WLBXpPGvvv+yT4E/VVorH
Ua5K5SHE6vSiyvbT8SFeTwWSPy+a+oi3DIT7KD5/HMjHhYfNiCpSfPOw18WuwHTz
RTTezHb7EF07TO8LB8nFjElT2KVZHEwqlDgQ36Owt+kJ9V7GgI91bu8800nqG+2X
VwDzS8YctCwEWblFZDfShyuV+wuAHBgsxvT2o0GMwvmqH2X16wpYxcR8p0rlB41q
veVW6V4SmH5lM0WFv1UHFr3fV5YYZvBZmZr0EF2m1HXNMYosj45tRJWnwfIhkgs7
KXFWxrw+i292npo/6maTq7/jpcFwUAbBw6fukdeiBQWwcDPGc71V7l14qJIPej1l
A2ibuoitI2JKiY77OPctUzpYM1zLCYGoOF1Sb8zWtVyNo76axvB9Nq1TH5SOpVet
VuVedaTGbS+ntFyE9z3mzTeMrlL9XhD2mZz9Tw6DgcVutcO+FHO+FBBZBoAU5toq
QsreavH7Q85dNoKVTpL3Zu51txuUfxrVJKTWrrnKv0vm+BYTvNrCUgJeTD+hsV8Q
QLhqq3wOa0w8EnfW3nK2C+wJCgt3/DlRoHW4XUPTVCqmDNUC0WQ1iEI+SmPNVuh7
ABBMTm4/2XhqzrpXbP6cRecEOkyPKixS+da0Qe8Atx+3bWI/ULAC6waRJs5iDU1F
1qlIkU+RCEtuXNMrDTwKTRkNNnL+Ea0oE5Yt8D/EkDOChXpFAKuhOvJxw5LHyLSJ
WGN9boEjKg9PGnu1sKCN3pe2XDW7mJcPHozyIZdQ/WrcAvSjRCM4yjxSX7E6hruW
GxjfW6ECLRlDaQLbe7DzjORDKYybnt8G7r0zQP3wdX2lEYPKiEK7a022CWIl5vsg
Wh7ugWqyUEeLL9ag+nCXlOfx0aE1P1mIwCiDY5X+qPbI5aCPwjRZPoYbRk9Tv9Fd
lOdOhrR3Nc295Qn0/I6GMKCPuuXSPGZMuWqiCIA1QxaYzjczFCpA+As/9qan1AVd
iaaqxnUow0KxkuNcZtJPZkwglDooTVOMhk/p3smkauNH4Xs+9sKEWSNIC2R8H3Ib
03fBVS7CLY8elapZVqmxmq2AQ+5nNbS7NXNmxbEaR0V9O4D7D8a2toOjE3cth9N6
xHoMYNzZKsD098BvjRV5y8dbBR4CEAmWPMjwfswcDV1uPQHAwS6ixxdxLQgubu23
3q2zl5TdjEmWI5IO8/pRsATUxYsK2Nw0usqasyggQ/8uIZNPpsTuJ8Ul6yCAQ3N/
aOsUMky1a+lNTCzYr8LtIxdq+zs1354bE55iDeSSo+Bt9WzvfQt/elXBB+t0gDtK
khNaqJebpwLbNiWWzc0/aIpPsh8snA9ZqK41Nbcwfbvhk3v7a5TgBfI89bQB6yXA
65t9CL7Ww25VDMAZB7q+hkYRRCR4KmxgCWSUvOxfHBOKHIDPe/o0u8jxVEi4wIKp
doWap/ndFFldm/2v3PjOJh2uuBoUILJnojWyLnOG2MUd8H9otsokmas1e9atHvZI
9yVx2yfDtRDlSuN1quH8DJO8hMIKxLEDY0LaS4EFd7Yjgng8pQx+kCuxjpPNBrkF
np0QT0JVfltr5K8Wr/QkgoRe6a9YXJyV8fmHaJY6mIHO+8s3cp13cJaWUU1MLbc6
iBdqTzejTzdoqaykKmeiH3GDexUbtfKGcWkvNWS0LxwI4+1JPtwuBbCR7w3wxXN0
uRxB0x5NqbO/Z76jTwuK8URXsjlBgXnKJl5SjZcgaUHUerZr0Feg/UzZtJO9hTFn
j3N0A61AxiRwIlJcES479A==
`pragma protect end_protected

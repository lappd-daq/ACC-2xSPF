// Copyright (C) 2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std
// ALTERA_TIMESTAMP:Thu Sep 13 06:32:40 PDT 2018
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
ZvToz8TpVcrZelbCmGdTLuX5fhm0GOe4wBC0QIf6v2xPDYIXyeX04iJtZBTfgAFF
lFj/H54208JxJBVLJKWlVmD9NJNzlk5Bxg5y4kBCFWw8kJQsfbgmbQaelbh0Q6wG
3gqKS+f3mnY/owinx6jBNglcMixsLF/nMvJuMAVqCPY=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 13344)
d17DH/YBy6E6eeVEux5z02BRbayjTGOHslBVW09gyL0e/5RpwlGQqGGUgKBppihL
vGtf099neseuNXVcpjyfWGtjP9l5SQhP2FD1MA37Nb3ZFXOrtISa+kUTLlaNblI9
QaFNae5ewxwaftQMPH3/bh+tmeED+T7mPxfKfezI93h3YrxxRMKTn/9ppj0T4VUX
b524CtZRdO8yFBOGAehF+2O1SjY8F0wf6PnKena7e/EZvb7Nz6P7QQYewOu5HwPw
peksTpvnRmZ3WPQByaLLeF6lLyubp5LouSDiV54xVVNsuFRoAP7bGVziKYvZ+jeb
cwg/e7C2l0JPSatNN8EHZpKJJ+gf9WlknR+McrFIPwfJgBDWbpo4Ll2DdCw2BTqo
cRkOb2o6Q25DqvAFNS3ycP+42Z2oZLB8o4L6njn5e8t99omAeNJkU+QovQSqZltK
ZpQ9CUjUHjLJy1z+EqD2nWtoHwaiIJb8mcHFea3+bEUiVwezkZ5MOu4hYK/N2hww
PT1wSulvTm3lI8wPRLiI4ExBHnTEhqZZ/Zuk2L/sI0TCV8FV6U+8pBUx9GwAeX+j
jNc75TB50u3UhHasqiarkqKeYf0/gavaTdnutyqMLjtmask8P1H4apxm9LeLR/m0
Rqo4Wun2e7DPPS6jRDofuxeTsg56vdTo7Y+M+UUNd22NvAQqSPgjTQzTZAfoHYHV
qNiYI/AiswBSKoGCYTECiz8sokir6P8csnAQC1bUcVHNl7DQaZRNQzUGYyGJWmiT
JXUs0pAsjfX0niMrbxyAxu/jUu7gA+RtWt1dqYo6G0ujpW1Rpz01A6qGhCXwBxBB
n0qs5yX27ZcGIkX+eIC6d9GzWx7b3OEUHsmNeKBEo3nl4t8Z8hvcy19dedGU/akP
OBPKonvcWC1V56COO7yeC6kFBB3PWyd/D4jl71ZvY211+OhyXvqpVevNkWarWJY6
BXuePIcOcboQyweS9H1Qtqcvmaz+62bmiqMv61YSZFmhBpT0QXKEgs3mFLAPYF+X
XKOFWexm3i2BN7r8KbRCc8KeZr/WYlEDYQhCEhfXr8UeSxoydF202Ev2NkSgbOZd
5j+UaZHciyS+ZuBE9DJWae/4Vzz9qO8M1i6mdDTPww1I8QM9Vf2i/L9Fk+AD4Xvc
QxTURMnUFQxMadSpLepSYvc17wdPMfNhIv9W6oi4H4D57pfA6PKoz/sh956gXTbg
hQDKyPWobSBE2JTJxm+qz73P3t9PyzbdBWti/uTE6txq/iXr9mBQqnRwq8AIYibY
8DuM+xNUI8XAUldDo96h11rfrVk0Gf71EObhczUz5JyYvCQChRDz2g63p/9X+IBZ
oq9dNYvVfLE/JNFaWewBK/L9P0ABO77ST6T5mfp3d02WFQkf/ybCTprlr2e+ff6t
QRCvx010KxUW1U24pp3PJSDX/BWmI5b7Clgu8ybs5wMXa3/ZNrq7Z8CpGKN7YsSL
g5gvTmGtlcPpU9X13MJYGW7uqiTiHoBxthhMLpk5+BdPjTF0DDdCaBSW/pwX8jgK
4uVBe8Es9ri9WliYSu1fiHYBXvG2UALKEmHMpQ2hK0GvES2VGPMXv0Y6RsNcxJQz
mP3HktOTbZS19PTCUyVlqySU6ifpSvGVI0vOT/i3z3p4mbulnd73L2lv0+mrtcLL
0+zl8gGayS6aNcuJT7iReePkWVpTdMzkqrHX5TQfUQk3HubMK6GfzXBnGX6FcL2H
xNJ/0HyL3DRYcp6HbNsR280Cu6d4f4kdaBMhV1WymfFu03a9IkOjINvU+yFAvPWc
OSPbYx2/FMfBe2WU/vTtQNINGyeNKS279cSGDh1GSQlbrKX4EeyZQuK2+bZbpups
TpCGlD4Ixn6U/J4PJoFYLyf2ebA8AgVVu8A5srBGdCs4nqdgz5yfbV/9RouNrL9t
of9jZXjUYOw+TPSIzCgaAbX/J695FRa4vfKNBbGnFzlCMrF/tq12rEAKgrvOibVk
2y9a1NT3uRtgU6Og/pEf+BFwFjY3/D9hR02x+Oj5Of8Z3erFZuDhFq2FAgI5PaY0
lLan1mDg/eMjLpPBGGfjRkpRloCfTyxhbIuCpvuzPMvODc1NFcej4ahkcqSK8OoR
/O2TNmNWn6G6R73Nv1Wv76FSDMlm3BhAH+oliPTrR5k7Mev5U/7umIlmrRxwGoiv
KuWr+sUjhUlWlpv6/i444O+IAygekPbAKRMmSIp6buZSopheOuLZGqJpUNqRR9kJ
i6+o0eWDSFeCxf4QebGAPySlX6D0V7+ImQqGJE+sxOsz3y77fh3m45/muRSF8ogS
DM65E0gFVaieE+kAgQxN5tb+noxm7bJdiumrvy887Q19vMwzAm0x4hh4/t7b+rn4
gLjBFa2A+shUzAHkMwe/Oqrtai0wyJDANbl4+KT6/ISYzGxIPwL4otK0B1X3DpJI
X4fVPmY5R7whaAoTvHSkpS6JvIDl2J6ly2KfqhrMlmnZn5FEkA5xpWYKQsdhwxHQ
zcf/qf7psF5mTwojIMRZsekPjF1Vf5D3NGkzAcsL35BonLKhrAeZ+g20P2Hixyhm
F7+//jhvPZjYTguPi6d9DKs7BNR9bFD1MhTgW91158P9u7EDZxfmJQeP62pblJa8
iS1J+Pem/bp8hkCCWqqFLXl9WlFscKk3NAC8TLRQ+p417SkWGt0dcvf0MgCMsmrG
s+stdicIM8ZfQOYEy2U7aKOqS8sB1UUAUs6wsdYQdZ6z9jaYVdox9Zl4ts6SaOai
RnvN60FPqe2irv+06Ag1Ld6FLDtDPoNHPj+DUWiacL3WMSoxjwOWbbORQ0ZAWVVP
FoJrxtaesX81AzOVB8ZEOL4N4Leht7ltC1oLD70hEsvaNINQm8Nqgz7tENdFh4nv
lh+lC/+RekwjGCmwC34bAZ2ws79X9MUU1chhemu2lHtNAKYsBaqjuSR5bSzYx2RF
KzWNbO42xcC99Ihyg5OoIJwTBJGHIgOIH8FRiL+98/lk1gxsJEKQn5DYsJM1ec5p
JU48Wnewenx7bhT3Gog4zaPdSssj4mQ0mFYVgjf2vx7wUiZADddHGCl7DHL8jA5R
3kDnVKjpw2dOhSgVUTOHjdY1+vodezAMUr/UC6+RvDLAQIEH7DBu5obQTDz2MYFR
Upk8upcTbqEIC/pb4nhnVg65+mJJR9O3NtZPnbZPgk5+Teyv8WLJO60FgF9e2K0d
x5Zh/awMKCSjGT+gZYAqcalSWSWnYLxqBG5zvoHFz6mh/gOJE8Veq8lxQIMja4yh
m+d87U0EAivI/NJTSI626zz4freYh78ijJgBfoSZ24UkBOrhW/w0yjo4oLnACcbD
tFxyLAdQQctu4sGjkMJg9NE2M4ZsrWXnNNW2xfPvUFTiC2UVRqbs9b4O20hYUWjS
kNVlPrRtOGSLxufYHYjLnoFeAGjbT8eJkGxdg8cOe51ftkl8j13YSd4rwc+uN7fC
FpcmQa2B3hRUVzw82xXclIFdWekHHJp5DkUT+TRVHBAS42RJMjui6AaoRXbAZKjl
eLGhqdzDLWJQeafmVic8bNAyoej/a6aFLM0zVaG1lCuBptBKqOh5nzR2xLT5UlyO
TRWEtOvkMdng7AVR3wOSokIH/sWc7r/YXuIhvmVtccQuJCLYUZ8Eo2fg7Fqjqwdz
dPCJ2Z15JO/ef9fUtt21u8rVVk2gxteCIkaNZNTmegvywAtGKQOep1ZnoxVgKVcx
cfHPfkMiCXG+Ei6bVi3K6RlHi6jF9FN0HbyJoBcjFIqWfVrjfogGy/9e4bNj2t5I
+7a4y/lOKCP9/WHN/pFTJh/iPFMijvd/sgIJnK+gfghy6d3pWTCmW4GBJlmXtV7x
A4VGdL14z2U+qhyykzRR0VQOTiYVW03tNHL3kpDtck/AVlY/wBe4ZGhl6HZLqNSx
QHjGmotASoZIzD6/F3RaQk5pu9R4WalbnXB99Z5Du327MpbHj+RfyLWceBwtL9Cf
mZyixdL35/VQ2yOWxGPy/NruIOw5QrPAdUF3MNZEPLH7e3c5I49s8kGeiayQT6BI
KXK5UNLHSQ/0Z+nEUrQUOZJ4MT1coOstd7CIw0jLxDuxnAmnM2vr9D1gYBOfF6qb
I1tJk7CtNp9LBXinvEJBJNVT2YkOPQNuX/ICC2Pol8j0GmqldqPmRdgZTiu/f6yR
/0sjjJtBcaoQRz0HySLj83Uo6Qpxbq8YRtSdR2TCYfvGQSCCmbuLOLb/Kz0DAan1
6ZOtzzjiOacxOFavaGpQsz6nLI/1dE4TnVbujelRknw4PMcAQDGFddTDp2rueH7A
2djq3wet4OiGjkk3BhW6lbEHAMGBGwTQwDiUyLTTd/4JyRxHNabCCSiCZzUJLsmr
HmxN22HUMVmEJWmOxe9cwKcVh1kUXT+OrXceC91psuM3hVe9av7ws+wKXQIUX5q3
FF85lNFGsCOePHYIPBJxh3Tu2j/xi2BGWzcm7Vxz+chPnzdgmQeu3py/Wkn+J031
hFpDOp7K0I59YTEdoLWpuXvx/Z7NKNpk7CTAIhWeEKe4pt+v/jpMUSBxjfZL/AUL
SDmzhEkuBDfgoE8ju8r7Lp4bgkHNep6fNcmXJ+Js7cmWc0iewNBgpKmRrai4H7l8
YgpRflJ1gKVK1DNukNKjGPIVP0SsFfcN6v2UO+QftbBQ7fax9GPf0weal3tOZ6Mx
qtD13pvo0mlvOujbYt1n6ETum4CXVdNFjCzci4j/BuurldtUBEE8ZvMELzvb35k5
jymdZi40FL0qXkWdNBAjlD0YC4kpIyIxm4+Ahi1zJFqM6VzvD9OQKcE5LlXAeO4Y
w0uQcLcJMZZR2ueUqPv+2uWvItYnMaW24cfQ0iH5lOsrAc1pa1i+0AmLH+Ki5Izj
v8caVTJHbrpIgxt+otCLT5m1I63RzMOPwiD3ToN5MXsxTK2KJBURi3xWR7KQcw76
Q2yBlwnEq7BrjtFbfIfZo42Imex1qjul8beYmeLY7fFAA/6f7amvoiZVAZgjUiMr
042HyFPN7O49YKXotBnSwxvdLeBjL1MGBJScygwbtj4CNoiLqfe+n6t1jfGEOvoo
KMRknzqNDZ1mRhWXio7MNEA0buS0tO9FMBAlXo9rhFgmT8cGEurGmW8sA4AO23D3
1VAUm2ZLk2SnY/4vInjBwTTiUxvb1TX9deIrfyLZvYaGodeBZtWh4+OYH2KT97BT
u/H8U4q9mX/bTdo0QTkAuwezIY3tomHWT6ZITIpMHUMRjTcSkO6k2Om72lIoJT/t
2Zyk9vvbtunjDXP4sfzlFHBNs9DrPHsyQhwixHuiQ1qFJS1iIpN+H5MXN6LD/p2c
yLIQE9lL8hYbTGZlUggZ2sHu4609pyyHQ4Ntkg8rh+d+tBkDuV1uUd+8MJ+qZuDe
//TM2xRiqwRl7hzWmqSauVIOQRlE3BQoOYxgHZ6/8g+4d/q6m0eQu/QnNtHXH79F
KtRSJSOM+8eyxr0SVeqeORrhcFqk8p7mH4AHvaRklus5HIj+tVhiEFy/j7PDKpyG
04+ge2I4TjnDMYgwHhhK0xFQejaUT9foaDQbwnQtLNCbRvYZuLAn58KK4qoSeVNo
DArMAm8plC8AGo23FdBRlhwOtCerEKBaAIxakt5IB4sTdKhbOry0yShKUKzej/1D
Y5jIVuarwY4Ij1A1QVVvu+cqX4siZlvDdT5JIYsSu4SFfpIhMiJIBag0aaZWi7JI
no6AqBQ/fu9CCcuNelFhvcJ74/JeTiCfdg4UywUhPjcqUbvqyIf7a5IJB2byRVVD
+vRo64+RpKuQCU3hNSr+VFYGG3NTT+0t8tKUHi6gxCEeU/jkFVzwAy6cNKsHfOHx
40NNiIDSdZJnlgG/S17yXaiNcIBqj1D95WWVFvaPHzn8ttRzuJl9iBlbRGp1AJEf
U1lhgsH20FyZ3SOiWZKwP86YSB0GxQg+HBq0VGZTAp+x4WPRpfj8b6Ezr4eECUH3
oHVJlS4UQ+zcUMkpVXHbchcJAPwX+vJOBZLWIsdYUv+IXjlS+We05SYrNta24k5a
8RLrf+Jo6Ohs7LhhQlBZGFPwp6ijPFu9rQFDXLR3++MpBp2FZihqYNiW1JP2iGkz
zw5O2/oovHJrpT+JaQXXe01ay5Nl6i9E+Rxnp8hOJJe1nzAmPsGNl6iR9c/alj+x
QFTs8/UIKPt2fVzDntyuvRpUC436HExQvbYqW2vzqaAiV0acfVj++4fhYjvr5lZT
qCGEkQyHc51pNatFyDyLCxyJW9jEDbfDBw8D5tPcMe+LE4KiAE68guWntQTM+XXj
qxNo5BQU8iNSYqk7t+8aMEnBnAjek/bHDeDGqfNi16sNWJaPBU+Csmf2TCn5iHAi
wnSOJ5hmuXa1Zy+zaDT9ajtDbKwfJFn9V5o8T4tAiLJfuR1NJxaDNHD1+eCxAy+c
YXoR6L4DnZJ4gvOirn2WAK4mBJ6uQ76iXxOXve7akd4hHGjGXgdyPXbDA2LnKfVe
8fYlU0GZlfunOKOUZiweqktoBiAsANp4neBoc1ihs0NKgZXYsXuBIYdWgEAj0yn1
3GHocGs28frJXbNN9ICfdPvAPLlV0rMm2Qf1YkPK4Ns2q5K1Z7H0T9gWesqhZiSr
YrFZmTJ6IDBqCwv5pVrldNenOEozY9bK95c3cBIsx901EGiLwVyKKMguFnlcNuuZ
Dhbut8y1fCt1/hIsJIPx79Sn4Ni/ipUDqA/+uZ9UsZJWRsloRrGadyRAT73zdkMp
rnkPaTQSfD8W2mA6/UCu4x8Qxxg0cAjYaWTxjxSe2okhDdZz9J4rTTQWSo34wE9r
B2qBpkyhb5DpUEmbhtY2Ew1gWWCTjoTrLld6X8DOVVbxrZLf4PGoZ6NW3cyO9v53
F9U026OJ8H/AlxPeqfZNYg5OXjrh1nN2IcgMZCr+no1ezfI4VOKn+l4UIsu7GVwz
VsZvGLXi1N2zyQEt+kNaVNptSIWH67YkICzOHV5rnSmee0CLR+fTNaLUasWXCBiw
bqNh/b+aa0kfoEDnH8lBh3X+LDfP5oJBZs/yOaftG3y2l9JLX8CkLn9B/52fLQBR
cop541NSodPX+iPOB7VpyvuuIHU1ByHKc1b1L935UQrMRoXGDDYf5RcbPDmMcO5Z
/mfuTq9TDQuAtsaYOis75RUjIRPkKOHxyd0AL7+MjmDlim4wCPDJKxlhuu1R7Adz
P1U8ZtgNWpYVoDvQhSzoKzfVl1o0o+8gKXq5GdJJqo9cipJzcDw3hF7vZavi/fcm
No6T5BwEW65lFW+M2mYP7qL0DEgs2x/dCzLlwWVmfIEgRb/BSkvVZR12qzhP+6WU
85KyeQ5RbALLwY5sYvqexjoY3p3+7XMVs0bghj3eN9MPBaLtNFW/vqWZmOmJ4ZZ0
D6wD5IL3f1X4VYjvjCdJ0Yx78Wc3ckxoOI/XnshZwphEvPQJ41ee1CgfZYwAGkVe
B6K2y4DH3LizjnByIIya0TZTIqesuNmrTyeJL+5FCsQa6jw7BIU/FvGk6sPKPgyP
36QQhDakd5JK+M8/oRQDEMYeC60slQVinYf+pP+bzTAkY21/vewguwT/GeluWh7/
riE0NhrM6DAfMqn0tUEHsW8moAPHCysiU9mMXr9po/PUb3hv0zKZv7n21bquJSET
M14II4z2x0mynTKnaaq0LonvwgJ/yMrLwwVVwhMN2zUsPD3c8POFKOH0ZTCBT1gS
gCk1WaV5UX8iE2NcaMJnRnTsErwJTGtWSTcWRmn4kmaXxrjoIUSlhYUiZaV8uFGr
jnyO95z6TQ7qCK2CDHb7sLrWoCbOcyW4sRhCIlhflqsQxug/apZQBKDc+WPXm/of
qkrmIBPB7lrfkmo2rObfGk5ZbUua+enOl4jiUMEjqdn1RAdqoJcGF6inPwz1OExX
6VanquMkqZzFjHLOE9hF8dtDFvamrIs10CP1LeiZO7+zaWB9KrdtFj+Y6BELoqYf
BZPPjBZo28Yss/UWqCywNEm1N8xILuSpUmmHUWF/sy7QVBedvfloZFqKFQAqLh6P
gA3gdCZeufPF7K6LuGBDdJx31rxNx6gVaCpi5BehhTK4WfZ1HiYtq44js0VrjfXw
g2GYGkSzsWZUyEpdYGrA2fE1o9rlot8GwOMZCqkyniGrRH+sVKJIYctNGIoS75Qh
Wj4YjwH29QWWhMq5zm9W53xSVORf5tfSuRhzxyBjBdkQb72LkadMeW+7GfQ4FfBB
QNxaJZhhrSVfzIh8gpDmnRbCCBqXKP1l1+p3I8Vk7BwVrzNhK+09KnEKlYpdJRo2
maG2ttAG7j7T/jvxNR6bH3kCPHw+D3raefAQUlzs07Cxk70A81lpf+g/PQ+KeCnh
wEJmzPdw7b5BcYaMK3e/Cs6LrnS8l7aIZQYJm+EOgiMKcydGeMfjogXNbuiyOYSk
pjCgj4LfJSwjdXE0mVK5xXuGovHNWsIrJx4vmSyrs0io9l79mQnl84xlBZDYwRZu
DQiMq7BB5RaQ7cYet6PxzcyU9+CcMrg8loHRIBKRrNOU3y+wG3i5VlWF/rjjZfU/
GIa/kPpoWQUU5FDD0up3r/qoX/vsvwcY9i1AaRQg1kwawDwyCgBiL/IKk0i1Tmc3
Rl/HeXbY/a485/9XwKo9qk6GMo2h+zU/6VMDtT0dkmvcp6U5onihoKfhxmskEir6
KPthF3mYvKwBKV2yy7g6LiCM8hIasyAmsfIEE4yhCVoOCxT3zpdZJOJH0upu0HK1
7GHjkwbrc+XS5cXbiDqv3ONhrqmXdlVmzUFB/DN/DDyNTT0LDZOLPOunSkY8fXT6
30xuJFg3hN8hQ2Oyzo5P8bJgpOB+B9TebWHRxhBpGBt5EDdsxsXpRkUZy9blcvNv
js9qkoq1Eavtrq2d7L5yg6OQJpQjBBcM6y/l3K31fwX/lf5A6r7MbYvGFksWfJGj
Cj1V3DfR3UXYkCjwD+hzJzwwzooFd/rm1fdIlHRLp9m8hSGn+d6ASyTV/tse+HKb
XbEe2lt/Lhy4GK7nUie2p5mGb+ZfTXf5m/uSiMN7U/KVXHBAihgctD1I0uv4gHID
IfaOFfw0rNWB5h8g6noyM+gIymdnqpuIA7Vp9YsnvKtA5fZfQP1b6jiO9pWz2UNp
H2sIW/ANVuNlN7D0ZECnA/97Du9F9Iv44/MNI/Pp4uJfhS1EqrB2B8CMtNoNpKlO
v/1bTwr7kwC4RKxFf0PGHQikEAPxF0++Y+U6Z0/7f6cGPNGOXMDDnWR5Wnn71KH/
/PhdvHPtH+R9JG5eu84GD2Ckx43HyRvoo/1Su///JZf8Xpv041hZi4AcLMTZtlWF
SXOCuWcOdhq9RuGqJMvZtARiA3PjgXdmimx8Moc/6qv5S/2YClMoNnV1WYEJEtpq
pvw4urnnExSZSMNVBl0PWwaGbgo4yqSaGqbvxBXJpPKciIlEoWSdBrN+n0gd5Pgr
G2cmm0jKxwkZ0joYswr8Hxs8zcf7+V2oq1FgbE76+iVq/OwKRKKahxQofWuMpZ2Q
t+I2rslPHjgU7gU25rYMbTDCqErPX+Ga2Dg0ZoDnialWI/ltomAPjPrUFA0nsXk9
TX5IYe8NYdBQmbN+CgGIU/o6J2JgN80OdiW9nRIcZo1oIZyoo4UgVa8c8g6DtUrM
XfVVFPfoaGGUoMWVdRNqeVyWECcVC21LCS26g66GY/wj16hSVj62xXpG8rdE5e5A
orfscvH1pFwTAoJm3OQh9xItDHY+H8RpSTJoKZw3/ipcQ+NUJyosEVOV2121CHkC
z3s/WKr2STjLhe4DPSvKNrcv6HbG2fc3r4ma0y447gCgPvpLIcfM4ZkXQsbdFLZm
ATe6Y+j/HgjpgzsgqwevNwneweCjGcWR+/e4lpkpNnJD67RHYikzBh1QZlIMZBrY
4dtoWLkds5kQc9sZPATjqfo1eGbwMKnk837UtwAM/inXaJfHBgNzNLrLeaZzj1Kl
rW9wbGlMep+VysNSHKh+2047JYtCuP2Fd5motsoVeXvULrk8eLMRkFyB3TNjxFbt
BqwXKMPhZ5e3VpzPPplN8TLMBTU3q5B9eNIzu0TQJjjYajCU2n9S0P/qAzMDu7Fq
AlV+6IKHE54kDbmMxoQ9Be/NLwkZMlbEp0ME644b8aABlOr+O7/VYcp/VTbjIRZk
ylo1Pv/Vb2UNt7Un0BJN4PJmfy6DvlC4fqmEE4FZecNsvVkad0rQpR79hQNU/8nq
x5/Lr1U+XSrjERYwmpGlBuUlcUrRPMtk1QQ60mljzEBxJAy3qgTUcMgMi/+tkIWs
CEu26/SvI40Nmk1bFgd2fwXHgYhi65wWblc1HB2Vw6FNtki0GLZd67byoTFdk5Ii
dOjQNyoUBWA8aKu8BwgnhrOvWGDGCypdsg54D7RDCbcQbOJd6STRUC7zHvpWWfZl
4N8iDz57Zm0PjOg4JidTVhw3eQ6woL+ln+u8EtZjC8a7rfm12q7xctbVJF51bjUd
c59GS+tIzY2XuukFyCV4qWroBeTI5zrABSWdMHni3iVfo+reA1rbtyrjBYKtxduN
soVgW30QMMeLbWBUgYwwDV9baH7hVYiCTUDCJIZ+Jlz3icAA7R0/XBkS6J4ZSBB7
uMtljqI2NSzUuTP3PRbhiv83EN9hthDctA/W+09zWNwM3UCuo2VOX4+uO5ZDHGj+
0BY85xTdksJCGTiv1Y4iI9QHJlejBRPO2MMXbEH9qZuVm4Cyb2PwdPkaRy37ZrNO
4lOfWWapGh/XqjLZtFKDdSLX8tG8qJg17wA0dp4/KrAvOpATpHXTXiFZvBqPrwOi
npXwr2RU4YP22LusI2/vVdx3K28aYGs0LZrrQ+Ien6NnEhOwJ/nIJvHGMuzRbpe9
D+LJbuSDS08I5ORH/QnnTOLYWMV02LjdVesA+1i+4gJWRqbGp1o7VIdHm9YGIDYQ
76aJcv99Uky8q+tcaHPRzI4kwvOgF2QNgGSPXky/pdhARN2cEC11AQOs65rMYh0a
d9kUTLeRDuEZ/Ee9vK0ja6taLLvZH7zqh0ndcf4NtR/AnhfL7ZjdK0yMvqXOuMsk
nFXqzIvqmUisKHUiGKCxtkIOLJLpITqkJBoXpUiA8PTtk2L6eWnKl9K2LQEpuqna
FFFUW7wG0mDqOoweskrGQX3AlrEe0WulS8np84N9Gf/rDoGJ0WKUExZrm3aZPCyp
k4f3Uoy5f/uyGvp2OF5kN5Z4J0jmGKfLDOyd1DPBjmSLbNHSKXwQXARcDYyBl5Kz
U1eYtuvvdt8Rp8mvz0IEgvI+RMXbznnIBN/o1dYZixOV6ctDanLkQOpehUXalKju
2HTC07d5LEwGae2nHfJYu8ctILFhwapon1e9cO20KeCGg55u/BwcYet2KcjPaStz
aFLSg5vM/NNKt1bPspu0hfy/HObchxEzrIFy1yoEoRXwHnNmvvUN5qcVPu7JOIiV
I2XgF+7t9qf4TndWNmeYtmIeANhjBTzFxuO7bYuHcwQTJGkZdEMffvytrYsXIO28
OIWmOqUVaPr8POl25TzPThQwvdT+e2RrwmFu633oXxvvAzoRdOkb8lGrx5+7SikT
yeoR/MCXQkA5r3zF274eQV9wdtzwUoFYeLc6gvxT7zo+ZKXiSKKGCGMD7cNu/toS
bI/VJwYZfqmzxxi2WA/3dqBOTUmn5e3XGVpU7DJK4Rn/EVkmoPqsR1DfygmPQY2n
3xk3lzlK1J5BB6/txBm9/lJeTqxtejPNooHqZRhOca+/T/BwO62TR/jgYhwVuepp
qQnY9vqVLAstUbBpLugpXaz4kzxxC545ae1rdoLKWNv313cBMXBwCjZwxUPRl6sj
baurMFmm+wn4muGHWvC0Mdrjzyu0GFfhnvdvRvXvHq7mzNlN+yERPW2mTb+TD1IN
fVq6haJHaVpTuRwJ43KN5HvPw45JXJOsyiG7SOcLjzxzyClfRu2sqG4BtMO3UAw8
74DaM2ckmj/5Kvqe08NMQoyw98gdQcHswVBRJP5zvLhiZrtl2NVyLwGJooeAFN02
oZUp4aK2rwyfhr8UEpdeWiVAkjiYRMfFvxP9tqvp+CcvSVcqgzSLzidjQwqPRlid
nbQMMF2VEGXs+1LMtaPQumWvV3y8cuvDzWF5ZzzABe+Dhno0r8Gus4qycp+IDBvv
inBNfVg6avwLmBxGflmb5C2v0GXV7CFVDt83EJFcDfcIm4JkZlww6Fac3M7mkTjz
emmHLLMu8IAcBu2MVyVFuIyZ92WtzeFz8srjrK9H2IsnhX0QFYD1xncs2IoR7M7D
VO6rf7r0s72irmXIvqEVb8tNHh8ilo+pIym8A3bQn3PPCL2SIyfhsfnMiuwSTpRK
tnhQOTAWB0ZLuAAtp+IH0bvjkBdx+UHdSQtI15p8Bry0n9fq5f9PV/LfzKNWYJaE
FkU3E2WFwlL32i/uKbg+Q8kwA0GY5c12fTAbkbQe/GpY4Y7mVEaOusfnTkc5i7b5
wViwqb3bMu2ICQqxgNCZb6/WTtJpR6SHxgk7EWgNdMfxckS+n5d8Gjjc5bQKEBvw
aUbAvK34//t/KhFbXQdDsaXas5YK953v3r9FZja0vJ+QOP/h7Zn0vF+DfQKmqSmd
FPiZSnmp5zDLGEKmwISHL2Tqa/tUBlPcZUgcBYAeVVjWDPthSuhgrLjpyWfUcJFO
tsUNTVvTftmVKeEcs6URyxarSZQ8591HqWN3K4YZZTVF5npW/ZL+08Oi0EJGrE5M
oswgtcZP5LcZfXN0c9alrCroXEYJJHY8rP3NQhvJdxcXQCAy6NOoKnGa6y/jnR1S
2U14Ao/pViIMgciq9q8K1t1UZUCB15LPHFLHsPx5BqWgfDwd48CibhDqnWEjD+8L
oe9+BXll1ui8SgmoHxtmduV/d4p5W0/UzL7GlvwRB6ggJy71b6mCRbsEhfp9RZ3C
cKSnUxhXtnwkuIwP1yXWgxGBxRCNEy4xIHQLEIAbz3c5j5mJeq5hPnXzl1o/IxsC
PcEv22iy87gyxoLSaSes8I+Wf2NLMiFWxgFbmigUXXCGW9LrOWSYzyG5CfmvMzb1
+LA5w/j0vrweUAFs3tXbLFHWND1be0Z+9xZXP5mu9ZRtqQDX2JTAxvUUaNeJ3bDO
1v6jbZafOhK8JGloDMMh9zlYl/ELsXZFQVsMzR+8CdF6ZSN21L/SeRouV34YUcBx
/sQt6IwAxh7zoPBYMwtxhlav6udUeuTUs6g9PT0tQoDmPM3vaTylwVQYuJWGVjZ5
GxMze5lnL1oWIoxmwrVKPCTnHYhT/g3TKH3wJ4Ymz8c7JU1fNx51eJAZxgHRCfhv
oSRC+Pwp5C8+DwLNqhH+1l1FlET34djFT/3JbqnVOTphMtChm4FVmuyRJApTHwHd
VOmOszHfNwhPPCFT/IPI+y6vl59sVZeTb3OvU96F4QdWFMl7Kr9zgwCtS4s7G2Yq
9tKBEQJ7/SL3VIKitU2K5ukuDC3iUSn86Q44tz8GZnDXph9kOOUYu0CCAcbg6mbc
8y9bcF32sZsjK45lUqcXgpIt2AkBOx99Ha6zwo/C0yQulSMUuuGvepNddhI5EsUu
Q8rAVYJovH81xAcxTibTtTMYc28pVW/LTM+Ful1iBDf1k54p7bJoy/qF2QAxus/J
Lu2Ff1xEXv/4YkPgAHcE1FEpLORMFHNLgh/PPkmZOqjaSFAwJaZtNfDPy3d4GyYA
vcVsSdnjEVdR3OTcgESJnm5uhriFW0l5r5aBXgr87zq4vnjn9H+lbL6GZWZ0ROrX
hbiYztf6Lj2g7BCQbX2egCY/3hjkfLLx9YuDvchaNZykdXX8J7QPrivMKg71UJGk
YISDFLYjFuH7kR4xYnPGSPxG8POVP3AXpQINc1yXKJe8m9N6jk4LAHRCB6eGB4G6
k2UYpYdJu9C4IF3bU9Dl7+iqJB47pG4vLN3FJLFpbBnBrocS2+a0BXOojCAtlLm7
NFc5fpiVlXmtjbwMQBlb9ezxvoghEcWE0xAnMN8upM7ev0FXHhpkAB0EUimViUcO
r/25qovr7SQT5cq8omxkyOKOemXwYIhaJewYh8+mRTGr0sbaQOQX0ehNl0+i9Zfo
AwVcPGks6bjlQMLcsDBr17dxBmkrfy9RKBnfA8pNGt8u06NCOTjsaA+SZv3e0AEv
UP2XfA6mWDVOsS0+ZbT5UNxpzAsqx+s01OD5/t01k1ZPvWFoY7zWA5n7Pmw5IfOT
rkb4GLthgIT01i0uuoCU4HHH9iwHi4dzidZKWhJA9iFFwvI0kzSB5KlezasuUexs
dvpObEdvRvUQQwObvWiD3IipweQhFVzuARegjR2MY5hF+lekHddxZglmlkejjtf1
C6Du57zTVxlyEMckkEsuDxFPYalrPKAVcCbHCo385326ysJzfvP9Fp8+HcRYaXsJ
k+eiWb6YCyo60HJjGXaBHuc33zUi6tKnS9johMUhBvrTgSmNvpnkUAFBhvEnoGOK
/4iBHs+kaYiMiBtY3/+Hqw3e3vaza/MWAtue/hlUJtiM3FEDo+IaFIosH7K+2cj8
/VERO/V2IrJZVHs89qdQ1SiGVdi1ADZ7uXkHs9Q9qgnHkO4yFWpCEGlPPwCoH0ya
+/eQBYIWluPM/4z/xQQmqo6ITIebkl3sBvi83qA2t5P2vEY27cQBdbyRUI6hytDs
9dw90KrUIqmPAyBZesUSQuraWRTTGUqX8t4q8AsAzKBF3P2btuPW8++hidmihl+f
EFQ37FucQwG3/6d9N6N+kJ/MoCd/QKjU2d6rgiY54kxgSwyZkprmEynebbaIJe5n
XmwJrwWocvc9vVxsmU7x4I/9R03okOWzUroINpnpSRz5yetHCCa4kH8iGl8xV5pC
H155TYkXaZskTCP/mElpq5KvGzMhvfOFV8FTTsKnXRU4BQ6Iwi6pgrGOyrbIqgXL
7WBUdAaPEfGTYxijL0vY9PXHO70ohyBLTXPwXSGAkq9DM0+VbrXGHkRtdujQMfEc
0R+QmZ8Nv5vK9orL/H1jZ5tBpLJQj1vxV4cfilvw2oFEngYO8CBC7rcCH/YZ5Q4d
sFEyqG0zX6s1bF9nR0ES+6Twm3QcQgHhCIzp6bjfThdpO12zIfRZUKFnesPKMTe4
d+vTUVB6BN3IaBk6fbVyaqWA3i/OI5GJ1+JrLsKkHU69GuTeDznEdpupVpu/ADM0
ayjdgzK15GIsIyX9qcfuuJ2ox2QdmE+a3MJ4zXIwsQMWYd9ErG5nIBXJlrTx/ewc
kIBfuGY/tXclHOcj1+oKEHhJUSUnTh/UUMVNXZV8H5c8Nb7TjR2aduThYz3Y7kFp
vPlp73mNSF17LPuGfXGwNptWubiDwJxhu1ikq7KCSvBdIxTzxIpiZlYUWu+6KRDK
plc0Dk5EL+RuXeA5gimjjkGuvfVnYtzoYBD8lD2LKtu65NtXqztJV/uNbNNN8It/
QWZR8vE/vmwfsrnoB2ScI4c8D/Q37ijgdL8Uh+3xyWHRG/Eobwm+ZI31d5c2Msg8
W1VJQAYK7drOdGrrI0Oe9kb/jVKfPR0AvoZ9hNKBEz6dPAl+KyWBfWOxhd6HyHQK
2fPehF2DtzOHLc8xW2wxE8qenbVw0MBldsck1da/mRxvUoJTcvLxw9lOD6iH2dfi
rAA6jO4TIhiO9oAALcJDCZeyNboYP6rwNmIY0YIgLTE1R5J1ec8ygx+iBcZT57oG
S6wgnXMLLyuokvf44oOIscusya5tv/WSYz3Pp2K5WSTBpeOpJfYPn1DjpB4FExAn
jmGhn4Wtx7BRVwPF+4CKqw58n3U87xOVf/+GORM94BIj8K2dSXLwXf5GjqVXrFo/
2UO4SSyluErsyo9PqRLKJE94hVMHUeJyoJZZvNbcVT+bHtDR5BY4ziUt19lrou1+
92TEzLEW12wZesrDkbRcYKkjpDtAsXVPnio2RTWOdrerhoYHJoL6wYxiz+OjUXZZ
OYKjNsGriH9Cge1CXxzlnWv4wiYeYvyl7tqRKeYPk+iesThaA89IgITVLZsx5v/B
RkxuE63ToSQPXOK0+pfMQVRNHESOB+VU1OHH6yexV8sBrmPgAGJoc9zRqJeYPWLk
EriISpvPswREvlgwXbIf3B/Fya0MxKzeYJ+lbXBJwRPS1H8jKLJNND2ZIhJ32tAH
hZMDRnNq2dflC3KzlKttcNRKPet/1bFJgPe9y4gd4MN33GWtBCjdGTNxvW06DSWp
gtSPuoPB1PtsVokylHj2y8S3FgrnlfAGIg4ucTSb74BgQl0YgBOMfZhppQNZaH0/
UzqDnKyyFbnUW9ljO4rltrCzLKzIM9dOC2YkJT1+9uyBz/8S0Z3sQF2qdnPrtHLy
M6PxbZrqWuu+YJbza6RhfuVKjdooBWSSv+9xXi1sz79g4pxDbMtuC/vnoEcCWNaX
TQPbwBoE77oUc1MBx/lAr8IMrUwRoEcpkY3dMvFlcfynUC756JH76/w9m1RKYW3P
/qVsAV2P1GciPSj+zmf9988vq1cvGApODuJJi+c6kSyUE1M8bnZu4S6kjKp5FA/W
jCkYcEa4sxs0yDtGDXri5fnqJbI4EGnEz5mq5U6XMvoCbIvHU957/1kECIc6GhqA
YoPd7SoTm2s55purMJ1JHsc1wE6TsVBz4kdPoe8Rg+B+4nrPpq3q1WX2Vu6Z/E91
oOKngHdr57m61af+TglctzaYpEf11dNY/MraERQ8cQ9m0+9prCNImF+9qVMvNMx3
T5WV79fjKx3LfDLsKVaL82NeKG62jSgxBgtDiUU1l2JFJ6wOqTjAeqzpIaEe4NnU
yop1cTAFo4QjAwu28Oa8kRFvPfEvtA8a9dzv1/W/w9QqHFMLXye9puO47CoCr+m6
oUvXSfGkaU1U5VM5H/Vh5lzzS1iDEkTVAy+GBew/xFIdUFUsVBO1aUqTwUw3GnD2
qwg7rbCIVxn8PTp/GCw/fLv/OVcJufwXRr+/iF70PpMcXbj/5pZGtTreZ8va2nke
t6yHhZdSP6yu6Z3rpHBKUOFD5ZpRkR3JhGnipGl2RSjNFU9fV0YjXnDQ7jVy9MBV
BNUK3IU04JVA3J7oqkIUSMzOD7C4GrUiikUkmZN5LJCKnHk3IvLg5EGqzmbigzlu
E1KWCqLvv7OEX9St5DWcLtNoJHtMl2YgZBt5I2y7dzfwK7QuUnrBrkAjtxaPaoUz
Qn9z9DukLtMx5FRJYlqRpYMMICrNtW3Z7sV9SVKBJ0nGEr8srbjbLDr3Ln0mu0I8
Qfgob0QMRGPuXXXdqiRFiQUN74d3TGs/q36JwZVhvja4pB4VSa/dK5/zvOXJAsMa
aVymnwXEA6FFi0T1/jNf68+7ArKkbkRvxyiVbQUYbrCWuFPyVHB1nfim6stGLiNn
i3gjAKFYxbxH86oQ27fR8637qbn5JXDb6+lER3MnDtIxaO/s2AHLQg//gujXWjfU
68IRGMZHUNPPXzDSNOxY5PS+DCfp0vCQXHH4KpaK79RkRyb/Vy2wrnTG+jlV/fBP
KCntepEzWbAppNbPidZO7UDnm7N7ZdQiMcWJx6+wwwwqaOoeb49uR0cuF4BnN8cI
kE8dmZfLjEZJWap8c9ojhXsrFuwrBMznkEUERoq+RRoKul2vdSpzzEzSaOxYiv4z
i5kDP02vAEDjECpM4Ul77j9XvxQFFDZMQxHsOS8H55FXEUOPkmRuLHecqT05SN0p
yE2uHQm51gTty1sePt2gLSo4XtMuDFOPgkMwt/iMFsLvOOgK/82SpfSic5zWd0xm
FDtaW/xe4RT+VE8M7lm32c/V94wzGQhCWRf2Zbg3cgyquC1Z4xqH9MkmHkb4GaWD
Tzw3h1ae4klc/8/FUHYCX6LgTWFZPTT/Kc+oovKZ71tVf6FHESTHnDosrLl3PbEO
`pragma protect end_protected

// Copyright (C) 2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std
// ALTERA_TIMESTAMP:Thu Sep 13 06:32:37 PDT 2018
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Ov6LjkOJWDzVDF1BNfPirU+FLCl4IbQkzYdTdU+ZoMHhSowCE06GiKebEkJmDTRP
3drbXaGLRDG1OVP9/+hhAzsHMGbJqZxH4rvzVdi5lSs/jxRsWUqPZxKNYF9UWFnk
oCb5XQA4t1TaWWgEsrWLhKhCRvihUsUijMtEES2jRP0=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5728)
6FDHj4nPUaR6XCO/+DzRWR6gdc3aYzKYDOHdgNLx2pcI4dKBWEYjs/iXjxjJ+Ken
7D8dzUWsWEBZHaoHCqbFWi8YXyuU0QGGBXduyoV3TCgn47/+S+crwGc93CEXv3rR
RNM7S9o4UcqOpszBfYZK3RCbdXN/XU13m2YDqbQKQFj9OkyJxqAMWOIPK9BgfLbA
BLeGeKHIACLo623XVgdfK71lyG8U5gydbval+aO3f4sJh2caWNb/zJwsEiKPz86p
Qobc/OHZEHt8cxzzfFdPma5zQRpPF1sQz6Dep7G5cJemomwFObbUKY2s7fYFdtwe
aUVYdoMZYzBxG4AntgS2b8b/8hl2zVnEv3hBxrbSuBV3P2bCqTsJYWiELuDoZrdK
0eIQgbFo1wl8affvM4GNvDJm4wcforjwuxRSZQZCS2VtwTLHRpSuXsHses2UJUe4
YbKVGKFPEoBCSCP86nuOeKEEHVaJtMQT2KiLQizznNzFHE1C08ghbfmh41txIcV9
TdgCNySBuAMxAQHdEarD8HGR+26iWGqab9laVudPVKZnz1iuebHj6mSl7I0/RYw3
IZogPoYraHFNtjwPrvNGm6xEj4KjT4afZfMKjwe1S5suhvFuOgSMAAUsnZrHnxnV
fgOMV9FItfRNBrV3mVNHrb+Nrm99xnVWYlNKqytPyOFmYfLio/Had/8zGEKQmp1e
Blh4HZRZiGovzEzZYGuK0LOfm1t5mtXmKY3Fk2cMIq/q56rlUNoYLVlqmzySckVs
S4XAsjJ3ag+SygMeK55VvcwIR8HbnomSZe7m3+q0taNfFOH9K/erubXtgMZ0xTwJ
nlXMmNo9iAQp7WKn4reUe8HtqDDgnt3LDpLs1xy9zr9AkiA87pn+hJnLKghK9mV4
VJf5xMkI32FBtUihufyQe8xBcpyTgtQGfSj8ynaeefdd7BnR5gM6St9gZnf13WE7
VBYT0hURCFUmeynmgnLAvDsMBfcXFIYKzSPzfA1Nv3Tg0zQJlsAU0A61GxqpaAZh
epgVa/Au7GWsu/RiyveIJ95UsWpc/3V4peBcrmqAfvNl+3RI/yxwYc854YG6DcfZ
FGQPloh3ykvWlMaxhBrmWGWFT6Wx+YzNWKla3FFfUHMmOgpO5QOK05hdxkeN2FPA
JqBoMAD2kxvVRSwk4VNRRJLtKgjFfAWbNT7ViCE651N578bcY5GmlDalEHKeGITB
TTPVwiuX7CgRFo4EsiyitdiwKE0+t6YtH/RNEDxkCu74NF/lOzgCXeViQd/Yid2Z
KsQnyeH9Ou3F3cQksxwby0K5vVNgkDD3I8kVDIguPy5b1sR6uE1BHnGmw9swBOBs
WrdIv/JUr6aTUfQ5syeNEsvqQP0TkdXNCZyvKuZM9YchdyzTo5KCBAjVMLCL1uTm
fzpc6WWL+UVk+ThqUecZojnLwMlp8n1RNzeZKnGjk2t0Hkxgqf+LQW8mJHBHs542
gQWUt2vv+9ijU48UyiytFmYZ1X7ZoVytk5ydxQjHlE9rJpdnljg0t91eYnbUqJL4
sCEUGFHxaq6rsGknmCkna4ie8Jco+JJYlSYy5MFzdkBHwIab5GqZISBb6G0jycSK
N5xWSWOoHbQLG49GkR3SOidrSCiFAKDrng7qaGsLcKjOy8asiygl8kyfxp8cWsRh
92iLoTiF+myhf/JX+ML4gcq7EiVPuBOLBJfBQ3lrgCAEJ+Ql55aPfuM8CrBnCZhW
MJMEFfWo4dbmmTpk63NO0Ci58NTgFlaGaODntpVBb5aShgqJlLer0/uRb2lvebVP
yvCRMmYFMqI7im5g2Xt7+tJ0nExAURgGFbCK4/SrWCsR6RS9pdjXQXyiIg4uGJU7
1rzyOzn+v6dPlNMtbq16DcWjMr19zxJaOjH64XoW4S93HkyRgG03ORt3kKPO4sRb
osDcPZu1nVPY03j2839h/Qp7zXrDEthgteIC3WpFn4bLZPPzHxCWKevOZDls+uMO
ELLHsMvrXuSONYZ/mxozKX1WidxtA8Vwc6J49NEerlXgdgTBerwzUkoH2w0GjlXP
R37VdEn2wO+YGB4Te4YVCf2pdJb5j9W88JfhKl7zBM2GQ0b9OKRdNWgTvwbsqWZq
ld1jQaigtb/fWhXsq6x+biPeVKAgKFMOP3v+o9pPF6piFfxA/zuXv7wjCy7cRmbL
56q+4Y+hmWUlI3iqRiP4gtF+BRYP9+KQjsoIFbsvyLr1+WmThZjJEhJf8S6zXY2G
Nyc9WgkvCHxETp7IhZRnWaQhVA0JcOo8zKKZdUJZHWBousv8ideEM0pZabLxWVUq
jvRNo/a9kawi37H1oN+RFz1HodVnxYJ+Xgd3mZ2Ghz1sS2VIxWyDuewYZHSMr+/J
Drxzo2JsamD5B5iNN/us4EJeUokhBcFnF2dDpSKatHTE2vcUL6hDEqy/eFSuoh8V
Sx/glRP2ZxZDt3Sz9kr9vb31ok/q4YgsfwL/l3qsvcup169kxlVaqSPYqr752l4q
itl2dSOBz2k4MDPA0x3WJq8FBnnCCIQn8U913hSKWoQdJTUYLI35td+JNUTIqTbx
OlNwt93MFiWmkBT2cu5twd5nUPw6l7vhsPT/wiN1vTo3mN3W8K4k8gHhUMtw8JAb
OYdBxfvz1DhgiPmXVPlUCRHfaN8kPF7WssWI1iYXut+rBBkMhUNQ+AQ+4NG5qqnp
GDWhegtNO/gLXG1HDx/XHsC6LyFhYsP0fZ3b9+j97dzcIQ8dxhfPE1dP55ahJSbB
L+3OZuF2WJVENsqG12DePl5eaJJTg13zPJXocqU+EpODrsG0EzYvEVGKDZ3CNVbn
HN85mTQ/WmgR7Dg04fV+MjRhmE6rYtjU2qQgzUTD/+D2ZJr520+whqgGiFdFuX4G
R0R0/AuMX6xoSql/oC3h/nEuuHDGLGERpY/uwOsr294hT0pw2n+7Fl3GuXAhVlPU
Iuu6vt2/S38CKRl0d8kUKLxY12BsBhgqDIjSA5EZOXZUPkJrA1qokyuF0jQVAthi
BnddkmFwyqdzGjUtFVnGnU94aob1VMkLHN8TuV9r9g733UQg+2GIoHvCPmFt0m0N
48FcjR5Pa66U8228twURaOVC4y71f5Kd/FRDfo/C4++lPc4V6fxTzk8sjRHJsOoX
AOVR0zdDtt54EN3OJHpe17IWWk4MHNDzyQzVE5zWFNsZcuJnh5zeX2YvBPhxfoMt
Uguz6T0Uz1dQCrsoCr6D38xIcCzE402osCBr63VUyCnQ14nuVmQcfAqDEkpl/mhc
slnePoXEivgSptqNVZxuZsyZRvJO6GqUv+POnHB4DbmmvMUkoMSYUGCLJuWU+RDC
xO5mo8obmU/R4Zc2mzWS+szSo4CdmmVTJo8HLe649PFca4Jq43McYeoGQ6gokbSy
uDgcHt0NBD4awfczkn9RhrthKuBiM+T4kKCSvvEqX4U1odDurtvSkRtucelW5pVP
lIEpbWyB6LZ9wy+hWQI5UMh0xsFuCp105gYsDRw74aeeR+YABQrmw0GV8a+hruFE
sbxPtCKzqTJ6dJtbfyqx/IafqdEfl/Tzc9YOuoBwUcaEjASwKCeWell0ECWD4EIv
6QghO5uRj/ak/xfZr/j8SJDL2jUzQIZHOn0W3fySrMs07nvjo65LSb33JUphnzhL
SRqX3hDTVVCgnwIQoAjHPHXhb0YKZBSuFejh3cjlbz2KARF+FNECu+ONoz+BOjxH
RBNkGwipuR6DibcHQKtRidlE93mOs0J3pqHYcOGQR/5IzE2slzv4kZovcZRZC5zI
ItvKvLN+eWdHP0a4j8lOubVvQvDo2tS2w9rOFEDyjWGIU83P8Jf+YPUEe35ufJpK
TUhmDOPFwqP78unVEspDc0cgk/Lltk1wQsGCPdJCo4oSavV3DA0UWtn3TVBtOWVQ
IyQmmeKd6wY53nTsu8cTIkVJCmyvEMNaLo9hfHfOBZ1iqSGpQJG+qfFnPdAM8PB1
K5oa24EZ7kV3oNvyENBtK3jpPOLPkjDcMrKkqAzkuFGJEcA/Z1l8EzQKU7Y12aza
Ce5Q4yfgMFKRtMvvnk8JLADfOFJw7UrNvjcG3X9jWC5V8JdJCIcaNwj/KvF+fet8
Xl0eNXFSrIV09i+A9tqXBE1D7cPZruEPKz1j3+djhHPOjUTGFaaTyCGzm0IrGGvz
5Xfialw3rlA823AJjF3t3XDlvh21al7ko8mtk9Nu8a04cTIL5L3MSbz1BdNQVxOc
+nx+1WiKVIYh9p88zv95G9yUcfmIwkXnQaWIOYieUBc8+YfoShVaxkoxtKhsQtYp
wD0D1lMttQ/yvpdN5ocqHvAvulXC/L6GoC51ihBWFhSiI5EpQR7ECGNcZJQZ3NoX
GXlwPWBSFA7F+4n5RrmMf4lIeHpPGCT2738CBRuV++UL0DpnlBRRWZDQpWid7hcK
PgJi98pmVDOcBL24op9uXZhf08j5EnVBKS/Jf5C8G910tf4oTkwaxEZV/RltEiAH
c5AooFLqnLzEidEK0FpRrazZABWehwPFYJae8zCqErxDT2KEpJsx62Um/lyMNbXN
S8rfYDC7S8kPT8bcVWf8xdRIfHFmPJnpGLN3aQMioMIT6dkODYVydxVtWybtHZ+P
Wt1lDJW3eLbitTdLxwZAfgZ/rDA1GbeAZo9nGLO1Lc+z0CTi4aBgrs6YHtgVcgyB
AMqk1JIQPcK1fccPnIWdO+15NJSXxMn9bjx3kR3dV0UaHcAgmdwrVH2YKIJvzOVv
MBhY+jbu5wczM4s+oeWVRwl26X5glVfVXcdKhGt++FYSYZ0TElaqW5ujjqxPecVY
npbHZM8i7q8yFRu8KwzoKfGT/S6hUTFbGP5CT0cPc3eHshf23jk/aME6jJIX2D+E
A/l+Hh+S+H1AGriUIp/Gr6vocx5INVW2EEer1C0AK6nIFnd8jb56I5XVNVSUX2Wo
bNx4c0PDLdWhvNOFAdnxNsZTvVClEKWyOQ6RaO4+S8VVyoTZDuyHKy/9BUA8zGqb
Asg3/sVfvP2mX18MhZW4+rtfzVUhCm29+5JTkuC5IFoGp2y9Awjm/a6iQowRiob4
4jxGTwF1GNuuLeqee6k22jdJL2Js0mff7vDOInKv6omLLzCjzOA820IRxenwBWQo
jsY+8XJaxG5Hp6/e4eV+5EmeCZVgygTisschV8+OXWL5fIG9i2xPErXrVeH554Cs
ZmLZrhRAaGJtyZdCcvwifrjCWHB9ssEoLPchOP3xadYUVSM9kGqUrnBP7VxXB0so
0rMHWBgsJ8JBRn8e0kj30GvZP/yLcoRlGJI9hyr435hCaxDN0m6CTBApjlbuipyg
uLVMyESux57UmccbMFa32Yyweg73PWH/kaPjAW61H1IJpFyaqCX2ip3S6TFBK0SA
j9oqBrH+de90UM1d1wZfpOG2DbB6JIvzILHiRj+XKqzndhgzMFGUSym5SwQCVBuR
o08KA6iQUbVbS+/Yqto4U4wIqgsse5XNOAbDOg8KVlDqr0BMjdiEnDlOjlEAhwMR
Do75qQaz8IEjo5cLCWGx0s9kOjYghDwAD5+K/TwKDFDvCIFAbQf5rm5E6eDS2N0+
8oGLPMHi0m1GGZ4on9WgWv9rLy3Qt8WLbub3ItDKTfJACHnQKMQD8Rr4KQpbZ8+Y
CpG+Ash+5W4h2t0T2+UNmrWmE1zr3mbhccDOvWSJzmYo3rWbaVDpU4dXqh+5HMtU
Zf3HSd7oXk6B7KQe+SWxoErn8oZ/+cSlsypeGccv1kVfg/eFpNS+HvP0OliaeOh2
KLvdNkJoZC3eHlRxvieM7i6PFjlo77PChBu3XPGSshNTz6KBKK+uVzVgtu98fVYF
3jrXVmyWzMzRrHC5MpUKlLLJOks8XRqF176WHHT1X3bJaPvrHZU+uutISdK+y+pU
bs9CR/hfuDjIQDITfHWd5h1+rH8JpS/thEkVp5lXw1B2A5b+GAwYP+k+5O1NpPNN
N0058ma+0MgsQN9zo6RT2ODCHGdM5qbCyqFLsdleKw3QVpIOELvSNPSU+COb72G/
XaU7nAe2EfHcxR5hOMw+xHhjtG3tDt1lKlcAfrcqZ+dM+YzqQmdA+XYzVWpMOBOk
i9mUM4X1SuwDQqXQS4I5ZStRkBR9FQGQjs4oFDOqwqZ/HT0GOA9RJjUGs2mzgZ21
SnQL5m/c01EP6CpM8ek62FfP+r5VaCS+DgzgyIf8uoeF/91443w56zYa0r+WfCs4
g+/5kkjERVZLCmLEd/Plu3KRlrVLHuJATqFF/SNzxdgvcZsvhnnUb/Lm5DhoXd63
fJWrDManSq1htG2GNEwGyqcqXOkpt4+8IU0MNlNQCFl9oqtJuylf0zlTv4Pg0xPN
O4za9XZRkO8KmhS4rrWcZFpKPy+Oh1+I8rMEJcOBnfGoCFxCdpLX5hGc3JCyN+cs
wCDQKe3mXq/CUH6wnrs9n1WFnTaSIQjrxgZI5q2jiLrGbCCROjDxquq06DnmJnhj
oyml/Q2JRoUpEKc8khhvQdQApB9k0J05cITSRVVvRn6u7Ls2AwYIYjGu0xNDgXcL
1AFaQOKotONrORiL3mOA5/RnXZ0S/Ja0oB9IAkfsQT+MpB0DuIi455de2Zy/Zvbj
2mekDNCIdT61oV9oE05Iam0gdTdPezP9nRprq2CDa1Bo6br5oegyQzBEcJxMLDQd
HOFTHt/kq8Xw64cBwS2KlkugSDr/PXgClPof8eBfektdV3kFlgRs3EOE4dUNpxSy
+2O0qlPnCxFXscRWp+mG5/3fy9+6ttJylYwzsgqcXeP7wWPN2V3mRQQo8DCmWgtU
zSyj50C+pKK71JBL2Ws5Sm5hG1qKK+vHT3o+PorrExQBAA5Crkysdx2XAMYu/SrN
QXYBSJSWM4imfxyFzpe6L2mYkBq36krhPM3RI+HLXBBff5ZJwrHHgzJOWKWLG03W
dp0gHud09gf7foHHhUjIWVaFadBnGUbFvBNWZTueCtCsykeGhDHInfiuB3YrIYNI
P5gAL1XmwETJDhUPQDEsQaIgvfxOzy9+VJcCgpDCxVF6lm+ZtH1NvOzS48yQjgbP
oDDhDQLBWG296nFlzPu12XL4d28nIbD06l2Hm9SitRFSmiGKtl0w1oFYROXdjWyj
iyzO86Uvu0MbzHwS0hA3m3fwvtqzxgGVN83nEaaAbhYsdHLNFepJmkMzaeznxWY5
qNcwSmeqsEGQhmyuhPo1MTVCRP4ke1W343KQ7V+7E26QLYkwOVKuEFBKWoHQE9FB
cDSiWxH8OZqRzHHnIvIfn9IvSQK9V4lJoCOvXPoem20VwXiqPon1FB5vjAJtsGl/
vOlTDJpO8gxPyFxx+Z2xxiRrpV6rA6bJQd8safRh0qkzPXVto6TCDCV76V2dmVLu
H4p39PraVrNuF97qxXTxIIjinUL6/1VjQz/pxXUGx+tsH8v7gE7IyvjsU4D5uJJS
pinLiXGF85WkccvbrP8LFfUsB2L1D6nKvkZIMc1sO82j+ovgchUcmhoPOi67JsGi
PveKMCuZ8t9H4seGipFPbR0zBxnR5idtSZpv3+JzJ+Lnvb2O/CM+cdqf1z7mJODo
Vr7jaKHcTcfNpnYzx5bG9yLDB6cm/MpOZ5Z9ke2ZvBSO2zaB/hWSlmSITiNWJwJK
57Nl1mqsSxgIVCgJDW2xsA==
`pragma protect end_protected

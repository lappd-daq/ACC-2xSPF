// Copyright (C) 2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std
// ALTERA_TIMESTAMP:Thu Sep 13 06:32:45 PDT 2018
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
ibSg+AAN5skO+03dRq/YshMXgehLFGrxCwJqvPlRbc9k4zlDxNW4uga925KygUcn
vvSfs7pr6RqtdkNXa9x0K7Igb/eGeCYwpAGCUcRzAmZmOBwm/0VGkBBqBbIDABrs
vPO8mRzaV6448UgdeQxRmvOh6PpGMrImJwvMoBOJ7Ao=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5408)
WCiYhzzo7QEYASMhmbVMsnZFmXqL3DbuSPUmw1agMK5jOOHLEkj2hRJvGdqmbrHl
pmQiv/zHNGmESvSt2iH9fwfYvoqRzcUDNJHjazuwrv11u/1B0STNEAs1gZGRogor
/89Q0kXtQkV5bprTaML7jrdKzk7f/0srNL9UNkFc7rhxkx1sPfPLMuMaDA4WcrBS
uI7kAZUKRb/vgt+Xo+PyiPJ353A3RC6jh842uGpdUgOMuNCbsTjx6mUNGYVXgHle
/ILFL2q5x5J5EgtPOQav6qDPLBTI29TQINAnMIUZj7a3vJkP+wre5EliCeCeQJW0
+lk1vJn0y+Vzd4TZrcGcQ9R1RFIxN2bt7ZwedD3NAWpYSqbB9OpfiIlIsbCoziZC
eeAJ+btgdARKoldumROAKyprTZ1gFs2UczB/jW5vEbAEqj/I4WJrtD0ZSUcpRzSi
CnvSmXbEEP9Jv9kHOLfRbOuikPZ2h4EDvpO3+rrAX1QRK5n3AhQhyIsYV2w0rvG6
+f0LeuoGojdVKDYOzlRVklm4rjgnQpEYU6MGdl7g4xtOS9VBO+f380t+4wJ9xckZ
ygZ5xpCcMcrmrFG+ec+pSA9c2/jgAgKHga3GxPIbXem3VweGsRNFA5pqKjPyFHuL
XXmYwso++P/v9Zcru+JEltg2nrI3wkDn68+xssmSlLKHI1+YNR7RH7itt+g68NK4
SPeyIijaI6pHCu7+ukjEyEgJGJo7RbFNDFvxx6j3Ix25WV96CZ+Vf0pbLmka9cu5
3Khii/pi64sFH3yRIqWdIr1u9KvQ7vt2PytLMVP2hobCZb9+wfO4tLU32ZQGkYY5
onRpre07+nrHCsn6BPuMeaFgtY2T3Y0b9rLYt99Fqszilv+v4aVohJY/Vt/xjpbe
Z8IFi3pH9U1EdIXucvUn20kAHIZJjZa/wXikZe5V9qz5wSkV5hQetR+MSUx4d+mQ
B+0c0mTEEy4vYU52NuERvuEKEtCV0KWhVkwLscewUFLToOk8mLgfmLR8gqG1BLHW
1noCj6+6tOcF1kFKb5V+SdMKJfFRjKzSZpHAIH/zWYDoAYrE8wpVAG1GVR0pAKgL
2u5MYiIPH13l7qEMbg4XRJss387HrEkQTwm2uPQp87ZiNL3oBLMidbqNscw20cBn
+HRMKjYAXu8Gq0qqFz2f7Z9hNdbno2BLLtrzh4LKR4zjSWjmqw3+4cehmunc3873
bS9ARVzasEzgxGs4tCIwsLyseUDhMX3xtRcIXtiGddcPG6F9io1NFDJ2sEZr+WcN
Zj3NiuIQUmNi02RjnR1R5RG1fp5aWc4CRd51mft+riiABtXk/tndar3/QZgRU6kq
gZlnFLHaZazpcCK0Pz0/PsaYiDt8IrpTU/Zf5NAeeCU04/n6XW98pcrEmBT2YNpl
SpQZZewdpCNXQ9ivZwQZsW86xFthXUjl+SFsI5Yldi2ZF5HN/8I2AHai3ibGRvJY
htUQ9Qw104KVIL946cRJ5AW8g9cXZCy8WJihJ5kWflerZ9CdU8Au83pHd2+gRGlx
peAXSovwusRNftTSzuVOvMPo+SrOtNI5YOq1QUQoFgVlZiM/JnrOEVXeSluUgzu0
b+2xxLjpxk/E7BrkcW3c/cDpG20BbDBrUGvPS9U/76Hk2gytnku4qlh0zQhLCMKy
JQWE80vB3u2XoE91secdiRpiackixuidEy/2Hu6xFNJtvD5Ua6a2gv2O++kGAyZ0
82pLkoIndBA+zi/gvD043uAT+F4wPILa6i3HQKB9nFdvWexsZ8VM7JQ/E5RecJUA
9pI6a+h/GhZHeTv3oVCtVgv4tuCS5tVoqGRAoHuCiOonDIEJMYpGYmFfuTcED4VO
CdWp+wExamlT/9hk9ka9mtxRkLmgxkJfFoUByiiKJrtNq5B+bjfCoUCx/wX4qeJ2
QFSAmnu2R1oZUFGbcVNwOo1zxVNBQJSfpqzIfeBj1Op5UGyzWCBHECP5JERIgDLQ
PUJbWwNX/BFgucxP9CHfK+lG0FPAX6KxzXGWIuOkHGm7nwSVke6PfVcab8ISGzy1
a636XWkQkpXLw9thBnaZNFrIqmsZ0T1dvaym3T+SioPi2Nn1i3Hbh+BujalPesNF
pWdFr6mpkYZItigdP0sRYAhaEbtwJyrcrwVQ1w5cDauUdFPFUJY3OkkQjAwqqvqO
nq6Voo+4vYtVExH42dU0m3U8J0tt3GBmfNkPlij4mLoCCqYl2P1//qWec4vlVBBd
Uy7gq6VrSC3OpI8ZVCu8401KS9eOSP7tIS1QiBcRuII2auZjba9HuhVLrEyMTiY6
pfhdLmes+YE+T4CaTTEMAJDhHstF5GyIkDsbBm4uAOG+Cmq/5cswUFz8d3LkxQ/t
U3v6kd+s4m1sWSM8FwoSla/x3oYyz0RoEFPCXzmFb73fnw9LTiyhyCoA/FgG3EQv
6y6nBzKLru9tNU38oMve7MEPt3nvVUvGP6jeeR8GqKLbFZIUycUqvfjnSZv1Xk9X
COjqrVsNP8oS891B6U5zUWaK82BzheiVbOCS2oC7pAxtGQ0+1saT8XemuPeQk8DB
yd5nS6k7ggHpavBoBSzP/G8H4EKUtzbmtPgKnQMXZRJLlqTWhvK0PH74RjmS2tDq
KdO4mkN/ajGVPPv258WbDr6Z4ONGWpS8dY4VEmFAck5CyTAMbaNEtsGyX2rRjHJJ
IiWPrsALBh9/+p1giY+5EiyYcYfoXge3js9vW4xpRBEjLHDHFs6tl6SobqQ04UNv
BOQIpkUiqT7vtDLekiAdqzAHUYZKIZ6a9hgJ46hFDcl8HStGnNfZG6qBFtTwY0SX
HUSFeAEYZVbc6pFNWm1ynqqUg3iNdO1+UrcJqHV1homzDWuyVC4k+0EN97mAFpDB
Ch1MEnoyp5nGCwre78W26/IuToJBz17ySPs+rx3ufz9zj1tMBsfLv+5RhGdDiYnK
TzYBJ0tuv10Giox91v/9+7VCuyMTMEA+AORZYtNGb/JeAWuNpaBtMojI+tYCUaFk
2E9i1jqjLLQodNmWx10SVQ7TUxM7p4a2Ufcfc/pEjdByTsek4PhqXyc4nk4HuIII
1AnZWLvPDKrpx3gpPARWQ5WArMcseM6rPe5+dnsXa1KTSiVXrrKcnbfkIIKVnUtr
pWROMt72HLEd9nU7nHsv9bYuWxw04Gm118YsNwAEoBnYsEey09yxwOyv9jc/Fgi2
slEESea1vT/kRJh4MIh2vUa6xv5hquTau1QQsOhLCI/6lNcf/CDlhFrAMwP18K1y
tKGGyM83tPglNcvuJTs1iQdlr7NkYMR6L0B5sAI6JFH0lGiKj50PO8gj2F9VmvCC
HkfjC9Ehl1uvMZFHSyIEjitNoqjleQGwtOF3SYAsR1wG8n/DNT7U26ishANK008T
UR+wQdRQQXsXhxAB7jCSiXws6BWB0gf2+zhQza7X8rFp5anehdUdk5tcXoKo6YFS
9yussDgwtee9QqT5fqA79oHcakNPRxgwW6NjzhQ14BvBcynp7NWtuHefC6rVaq3D
WI4B9v4PxhW+8S110Kj9g0IHoAtyLqcY9vZTqnJtpR6yXtiSVle2/VBFz5Ew6RdR
/HFcozpiQrydCeCavQts1TELaLYd1592AF8slPXAWQLEPxo1fyTx/3crAeyj0Aa3
IlIu06mKiXt4wqTwx0JNZPbXE3h94i9sDDpjFuSRnC2y3SiJb32G8PZ9jkSnAA1P
Z1IEbrBjX/dP40zuhnRj8TRcGdaW+kw0ol5fYIOd4lC/WaMktiq+oZmni0JzlGFX
qm+UuQx4mYY/9eopZQ0YVlEYwH7ITEVpjKBVoglrnRgU/fUpRRlyMWnBdmj+a04z
Ciz5WNAQtDWTmIN2qC1ZI/Z+jtBu1GuEkVNTCkaR+vm1jOdOa+jnR6BpX0lqQ+gK
zeC4R9G/71ly1IRzFL3rIK7WahL8tT0utK5HiI7AVOiPsGCR4csejnCM9uw1cY0v
Fo7w7OAuNxnHSd9kTCPOrPfiGg3TSOx6bks3Sv07ipAKV5Gc00OJ6V9/3UmNn6ZH
6093tme6BLj0PprG9zHIT75LbmdF6H1BCu7DoEuDuVaulKkWrF7Mb9TatZcWIcqg
cd909OVy7n1OcWXZzXzZ6K1/II109jOmqVTW4l3v9Q9ycSuY3Zg7UAklufukltZ+
Tzcmbn287hGdtWZAMKMmITRlsExQzKLTHma7udDr4xHyAJNLuVVGEN23DZaBNC2Z
zrhrxzRCU2wDe9uSdpsGiNTOTwrGuKLjIJ1CIvCMKYHjiGSpN4tsDI1oe4pYfgzf
9Vk0AZXUMcfQDAIlrLaC5B1FisFK3+qiW4zCeeautc9JxP5/rkKDEez3kfyJAgSy
17kMFrAhhfmh5VmbivLmTCUab2IWqCZmzU/vW9Nv4AQlAIqCVjYmrHe/jm//qYBW
vItKAjO5plMk+7ayXXsGHG2uOi4FQ+DZhaMbusQl4X5kTKu6MCfPdiG/gimvPh52
W5ZVI6DsE26wQcNdKOArFqeDv4UJTUigZm+ULALph4SMIa1m0Yd7Iai1uGYtP+uo
tiHoxBn02FDK+DPaxieyWrMAVNVbxQslkTFevjxjuTpaIGAhAhrtKIkGPlF19EaX
amtUXGFAjzAgWrS0Qi/v7pfzeeExycQECFortURL7RYdy7ipKgQwDC+QHpiQqy62
5HHn0hGOz3XNmz8LPf/sZUO2GKPlt5/1cJ80XutjFVJaculSyw1Y0N4Z9XhOsMZE
ird+fM8+GtfhDzIWDxQfF2SFZqdv0FNY/9p/+ki+81XJWxOl4nI0KanTn203QxCL
6OvTnZz8KnTeYylb4MBIoe8UKj00BakQOuGVFo3iPaMm7QkXq86UlZkM4wR2IGM2
7FfsyfJH35tf4UstIi8qk1n6Th8hhXcDU9EzmKfEomVJ6vEWpKY8ZMUjH6MOruNE
ZX06Hige8duescwPTF9jbpIhG7V29NHXtEaZjrmtEM5HRyMrKJwr8sPWdK3YSBDb
esCvqLWz0mNL+iT2duG6mmFz6JKH+lqwjjkMhFcY+hofJ/jXwhPuteKaSnevWh4b
jEzfQdpIehDm8EnI1BiRqgHvIvXMo4yugp8CVRHYXfTy9YPnlOS4S9ycwk3HSG3f
0MgPwL4bLDLV17F8qrmLI0+4ejF+tozZc43PhugM8c1vY0eOIiVARIbCjmjKtXKL
9g6sFeUtcTRAcrPdnT1Af13OFO2DkrbMW4IDJ9hzRRpGnhnylia6zS0ii1LFHYTT
t4nzusCh4ZKfZlWYy/fjqTqxsU5y/jewkPk/ffFo8LI81QPbj4Ggxt9wG/B547BF
Dn14NzoMRAXYJFsQwXBfvDhzezY5O2x/m6/IZvsxPm+VvYbbyIfkDEhJN2mnNcv0
Y7fMJEqnSWxnQzR7ixBY8qfvyuR2xj2BL4NT8iKiSH1tZ22Gazo2EFfEQs2YXM6x
TdHs1kMvcr88H3XopNX7jKTm5FzQbj+2Ek/yEyCDoOnboJqWD6XzPNOerKmJSMHU
XCyBT4OSZC5/oJEoAtlBFSoM8AxEx78PZBKSA47nGjeUYtlUP0JH2WBPv11TUbB9
0SYUXAv6LeKOeuyFER4eVRCs9svaqtZohDBujS3UzMbXHNBqLgsD6FIBjdSYnTiu
wJej3PlqsIm8/XRKQR3XV98tw1YoCbD7D3/HSatcLL0agANXaKwWin8cmJU2+fAD
0c7zvkqNZ/0mn6bZ0mIWZ/3W4JjYO8aG8sKmSvMXjyscb0kLaF4Z+aF7ztuOr6M+
P0Z+G2tjLwW/MM/mAtEb00/Oierr+SSSTgcbdFd7XqU5H8bFmVobJ2bpUa1wIOo3
TX1fpQ0NewENGzS9NxRpcdmMR0n1kXAd2djFtW3x15Bf1hTKMj3zDdBJxFtCIa1R
H0OCji6ZsQDRung4vdfsZeaoBFowhtyVdbVC52K6VUHCVfpdK6jTNnxtuIoJkRjU
H0P2Dr/M/wRJqlONhVKATleL2OrIezqAI7B/TSHsBK/LQaU9+ysH3JZeFZYKa34I
7aUrufg0yInskIYsLkrD5YKRvPgIyIKtEl54u2BMc+U9Vvkq6oiyQUt1MnX4ZjNh
MDlNz+6C6RWYP88HmIqt0hair6a2J/Uu3GrnnmIjR3NP1pab62IFXuz/JTN3p3te
WeLHDfkiG12GL6aHPK8h8Dqbpt4cnZnbBbLUpAwgBZJO9urVBx9Vxknqhs85W9y5
4q00Lt7irXlCK0ohGLEbVBDTX0wAMLBeYsCK+dA+8dl/f2jrnst+2KZFs2PR2hsS
iBXeR8sZT9sepLR7RJOWI/j/5org8tQ52OSub9UPFu/D47+04g+XN7K4vN7XMQP3
LD03E/vmvclupbW7m06IQ9N3pOfT1bPMdZmfPLEX9WiSFUIHrMZfA1sWGEAwEvRL
PDtVUcZ/2110XNDgWqU5ldgheSUpz8AvKxF0q9qshjvNZyhK9zwx1T9JPE27T44K
Zx4xxbPkRplhV6Uq1mqzoBcKRaKMixQhEDC0uJE8fgiPY6LyeU8683Sf83rmxAR1
fd2Ns4KbMOy/GHJx3mB7+J1UXacAZtK+wwBJrkAuUK7qBoPvYSAMwwvDecnE/Svw
aLcXY+Jhd5+evxAn8bH4CKde25iN6vCiffsQRNcfNPrU4LgtAoOwxqa2BTh0HnVb
LtgD8ZZZTbA7O5PcOzGrYEXGHkWfigHLTUarrJRQDPLIFkfyLeLtnvqYpTaTKB3+
wpUA2vCtzHflwyYWu6ERhTvqvGNWV+qp+QrC4TOZspxZ/PwCQrye1tFk1nGhQQhd
8iKVQAo5F7wmW2atTecNezPwHY/td7bdSzbEhhcIBDMfueu3kP+6pLPMwhx5Zwdb
f1di9XQvZK+ARpsManorGpHmhj2PnBq/yn4PIzXh8ZjpovtAa54y+5rOf8EpbFQd
REzyXs1i46qx9BtzIFLHPfSAx9UfWrm8jQtqsPCFgLHbxN9N2hTkUYpMYWPkLw2j
F9d/IluCizlUBsJYkZh9fFfxp18Lxgy7YMF4pvKKISuqmGcikLLa6K7R1ASG+H8r
uSGhgXipGkz5cOvHpqHowngBn4O/GXJjWVjzj84EnSR31UAgm8ri+db60f8+CzFe
7Y/0gUMADZnJpU6b1dZC+eA+D+Azl5Pmi7Zo1nploeGFsFWmXf7nO8TAI8YxHluW
DuICD4U5L6vtHbndsz0ruEZiMknPPB1+1Xmgh5c+UJk=
`pragma protect end_protected


module lvds_rx_clockbuffer (
	inclk,
	outclk);	

	input		inclk;
	output		outclk;
endmodule
